module BPU(
  input         clock,
  input         reset,
  input         io_inst_packet_i_valid,
  input  [31:0] io_inst_packet_i_bits_data_0,
  input  [31:0] io_inst_packet_i_bits_data_1,
  input  [31:0] io_inst_packet_i_bits_data_2,
  input  [31:0] io_inst_packet_i_bits_data_3,
  input  [31:0] io_inst_packet_i_bits_data_4,
  input  [31:0] io_inst_packet_i_bits_data_5,
  input  [31:0] io_inst_packet_i_bits_data_6,
  input  [31:0] io_inst_packet_i_bits_data_7,
  input  [31:0] io_inst_packet_i_bits_addr,
  output        io_resp_o_valid,
  output [31:0] io_resp_o_bits_predict_addr,
  output        io_resp_o_bits_is_taken,
  output        io_resp_o_bits_take_delay,
  input         io_bpu_inst_packet_o_ready,
  output        io_bpu_inst_packet_o_valid,
  output [31:0] io_bpu_inst_packet_o_bits_data_0,
  output [31:0] io_bpu_inst_packet_o_bits_data_1,
  output [31:0] io_bpu_inst_packet_o_bits_data_2,
  output [31:0] io_bpu_inst_packet_o_bits_data_3,
  output [31:0] io_bpu_inst_packet_o_bits_data_4,
  output [31:0] io_bpu_inst_packet_o_bits_data_5,
  output [31:0] io_bpu_inst_packet_o_bits_data_6,
  output [31:0] io_bpu_inst_packet_o_bits_data_7,
  output [31:0] io_bpu_inst_packet_o_bits_addr,
  output [3:0]  io_bpu_inst_packet_o_bits_gh_backup,
  output        io_bpu_inst_packet_o_bits_valid_mask_0,
  output        io_bpu_inst_packet_o_bits_valid_mask_1,
  output        io_bpu_inst_packet_o_bits_valid_mask_2,
  output        io_bpu_inst_packet_o_bits_valid_mask_3,
  output        io_bpu_inst_packet_o_bits_valid_mask_4,
  output        io_bpu_inst_packet_o_bits_valid_mask_5,
  output        io_bpu_inst_packet_o_bits_valid_mask_6,
  output        io_bpu_inst_packet_o_bits_valid_mask_7,
  output        io_bpu_inst_packet_o_bits_predict_mask_0,
  output        io_bpu_inst_packet_o_bits_predict_mask_1,
  output        io_bpu_inst_packet_o_bits_predict_mask_2,
  output        io_bpu_inst_packet_o_bits_predict_mask_3,
  output        io_bpu_inst_packet_o_bits_predict_mask_4,
  output        io_bpu_inst_packet_o_bits_predict_mask_5,
  output        io_bpu_inst_packet_o_bits_predict_mask_6,
  output        io_bpu_inst_packet_o_bits_predict_mask_7,
  input         io_branch_info_i_valid,
  input  [31:0] io_branch_info_i_bits_inst_addr,
  input  [3:0]  io_branch_info_i_bits_gh_update,
  input         io_branch_info_i_bits_is_branch,
  input         io_branch_info_i_bits_is_taken,
  input         io_branch_info_i_bits_predict_miss,
  input         io_is_delay,
  input         io_need_flush,
  output [7:0]  io_bpu_debug_branch_mask,
  output [7:0]  io_bpu_debug_fetched_mask,
  output [7:0]  io_bpu_debug_predict_branch,
  output [31:0] io_bpu_debug_predict_addr,
  output        io_bpu_debug_is_taken,
  output        io_bpu_debug_take_delay,
  output [31:0] io_bpu_debug_inst_packet_0,
  output [31:0] io_bpu_debug_inst_packet_1,
  output [31:0] io_bpu_debug_inst_packet_2,
  output [31:0] io_bpu_debug_inst_packet_3,
  output [31:0] io_bpu_debug_inst_packet_4,
  output [31:0] io_bpu_debug_inst_packet_5,
  output [31:0] io_bpu_debug_inst_packet_6,
  output [31:0] io_bpu_debug_inst_packet_7
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
`endif // RANDOMIZE_REG_INIT
  reg [3:0] global_history; // @[Bpu.scala 73:31]
  reg [1:0] predictor_0; // @[Bpu.scala 74:31]
  reg [1:0] predictor_1; // @[Bpu.scala 74:31]
  reg [1:0] predictor_2; // @[Bpu.scala 74:31]
  reg [1:0] predictor_3; // @[Bpu.scala 74:31]
  reg [1:0] predictor_4; // @[Bpu.scala 74:31]
  reg [1:0] predictor_5; // @[Bpu.scala 74:31]
  reg [1:0] predictor_6; // @[Bpu.scala 74:31]
  reg [1:0] predictor_7; // @[Bpu.scala 74:31]
  reg [1:0] predictor_8; // @[Bpu.scala 74:31]
  reg [1:0] predictor_9; // @[Bpu.scala 74:31]
  reg [1:0] predictor_10; // @[Bpu.scala 74:31]
  reg [1:0] predictor_11; // @[Bpu.scala 74:31]
  reg [1:0] predictor_12; // @[Bpu.scala 74:31]
  reg [1:0] predictor_13; // @[Bpu.scala 74:31]
  reg [1:0] predictor_14; // @[Bpu.scala 74:31]
  reg [1:0] predictor_15; // @[Bpu.scala 74:31]
  reg [1:0] predictor_16; // @[Bpu.scala 74:31]
  reg [1:0] predictor_17; // @[Bpu.scala 74:31]
  reg [1:0] predictor_18; // @[Bpu.scala 74:31]
  reg [1:0] predictor_19; // @[Bpu.scala 74:31]
  reg [1:0] predictor_20; // @[Bpu.scala 74:31]
  reg [1:0] predictor_21; // @[Bpu.scala 74:31]
  reg [1:0] predictor_22; // @[Bpu.scala 74:31]
  reg [1:0] predictor_23; // @[Bpu.scala 74:31]
  reg [1:0] predictor_24; // @[Bpu.scala 74:31]
  reg [1:0] predictor_25; // @[Bpu.scala 74:31]
  reg [1:0] predictor_26; // @[Bpu.scala 74:31]
  reg [1:0] predictor_27; // @[Bpu.scala 74:31]
  reg [1:0] predictor_28; // @[Bpu.scala 74:31]
  reg [1:0] predictor_29; // @[Bpu.scala 74:31]
  reg [1:0] predictor_30; // @[Bpu.scala 74:31]
  reg [1:0] predictor_31; // @[Bpu.scala 74:31]
  reg [1:0] predictor_32; // @[Bpu.scala 74:31]
  reg [1:0] predictor_33; // @[Bpu.scala 74:31]
  reg [1:0] predictor_34; // @[Bpu.scala 74:31]
  reg [1:0] predictor_35; // @[Bpu.scala 74:31]
  reg [1:0] predictor_36; // @[Bpu.scala 74:31]
  reg [1:0] predictor_37; // @[Bpu.scala 74:31]
  reg [1:0] predictor_38; // @[Bpu.scala 74:31]
  reg [1:0] predictor_39; // @[Bpu.scala 74:31]
  reg [1:0] predictor_40; // @[Bpu.scala 74:31]
  reg [1:0] predictor_41; // @[Bpu.scala 74:31]
  reg [1:0] predictor_42; // @[Bpu.scala 74:31]
  reg [1:0] predictor_43; // @[Bpu.scala 74:31]
  reg [1:0] predictor_44; // @[Bpu.scala 74:31]
  reg [1:0] predictor_45; // @[Bpu.scala 74:31]
  reg [1:0] predictor_46; // @[Bpu.scala 74:31]
  reg [1:0] predictor_47; // @[Bpu.scala 74:31]
  reg [1:0] predictor_48; // @[Bpu.scala 74:31]
  reg [1:0] predictor_49; // @[Bpu.scala 74:31]
  reg [1:0] predictor_50; // @[Bpu.scala 74:31]
  reg [1:0] predictor_51; // @[Bpu.scala 74:31]
  reg [1:0] predictor_52; // @[Bpu.scala 74:31]
  reg [1:0] predictor_53; // @[Bpu.scala 74:31]
  reg [1:0] predictor_54; // @[Bpu.scala 74:31]
  reg [1:0] predictor_55; // @[Bpu.scala 74:31]
  reg [1:0] predictor_56; // @[Bpu.scala 74:31]
  reg [1:0] predictor_57; // @[Bpu.scala 74:31]
  reg [1:0] predictor_58; // @[Bpu.scala 74:31]
  reg [1:0] predictor_59; // @[Bpu.scala 74:31]
  reg [1:0] predictor_60; // @[Bpu.scala 74:31]
  reg [1:0] predictor_61; // @[Bpu.scala 74:31]
  reg [1:0] predictor_62; // @[Bpu.scala 74:31]
  reg [1:0] predictor_63; // @[Bpu.scala 74:31]
  reg [1:0] predictor_64; // @[Bpu.scala 74:31]
  reg [1:0] predictor_65; // @[Bpu.scala 74:31]
  reg [1:0] predictor_66; // @[Bpu.scala 74:31]
  reg [1:0] predictor_67; // @[Bpu.scala 74:31]
  reg [1:0] predictor_68; // @[Bpu.scala 74:31]
  reg [1:0] predictor_69; // @[Bpu.scala 74:31]
  reg [1:0] predictor_70; // @[Bpu.scala 74:31]
  reg [1:0] predictor_71; // @[Bpu.scala 74:31]
  reg [1:0] predictor_72; // @[Bpu.scala 74:31]
  reg [1:0] predictor_73; // @[Bpu.scala 74:31]
  reg [1:0] predictor_74; // @[Bpu.scala 74:31]
  reg [1:0] predictor_75; // @[Bpu.scala 74:31]
  reg [1:0] predictor_76; // @[Bpu.scala 74:31]
  reg [1:0] predictor_77; // @[Bpu.scala 74:31]
  reg [1:0] predictor_78; // @[Bpu.scala 74:31]
  reg [1:0] predictor_79; // @[Bpu.scala 74:31]
  reg [1:0] predictor_80; // @[Bpu.scala 74:31]
  reg [1:0] predictor_81; // @[Bpu.scala 74:31]
  reg [1:0] predictor_82; // @[Bpu.scala 74:31]
  reg [1:0] predictor_83; // @[Bpu.scala 74:31]
  reg [1:0] predictor_84; // @[Bpu.scala 74:31]
  reg [1:0] predictor_85; // @[Bpu.scala 74:31]
  reg [1:0] predictor_86; // @[Bpu.scala 74:31]
  reg [1:0] predictor_87; // @[Bpu.scala 74:31]
  reg [1:0] predictor_88; // @[Bpu.scala 74:31]
  reg [1:0] predictor_89; // @[Bpu.scala 74:31]
  reg [1:0] predictor_90; // @[Bpu.scala 74:31]
  reg [1:0] predictor_91; // @[Bpu.scala 74:31]
  reg [1:0] predictor_92; // @[Bpu.scala 74:31]
  reg [1:0] predictor_93; // @[Bpu.scala 74:31]
  reg [1:0] predictor_94; // @[Bpu.scala 74:31]
  reg [1:0] predictor_95; // @[Bpu.scala 74:31]
  reg [1:0] predictor_96; // @[Bpu.scala 74:31]
  reg [1:0] predictor_97; // @[Bpu.scala 74:31]
  reg [1:0] predictor_98; // @[Bpu.scala 74:31]
  reg [1:0] predictor_99; // @[Bpu.scala 74:31]
  reg [1:0] predictor_100; // @[Bpu.scala 74:31]
  reg [1:0] predictor_101; // @[Bpu.scala 74:31]
  reg [1:0] predictor_102; // @[Bpu.scala 74:31]
  reg [1:0] predictor_103; // @[Bpu.scala 74:31]
  reg [1:0] predictor_104; // @[Bpu.scala 74:31]
  reg [1:0] predictor_105; // @[Bpu.scala 74:31]
  reg [1:0] predictor_106; // @[Bpu.scala 74:31]
  reg [1:0] predictor_107; // @[Bpu.scala 74:31]
  reg [1:0] predictor_108; // @[Bpu.scala 74:31]
  reg [1:0] predictor_109; // @[Bpu.scala 74:31]
  reg [1:0] predictor_110; // @[Bpu.scala 74:31]
  reg [1:0] predictor_111; // @[Bpu.scala 74:31]
  reg [1:0] predictor_112; // @[Bpu.scala 74:31]
  reg [1:0] predictor_113; // @[Bpu.scala 74:31]
  reg [1:0] predictor_114; // @[Bpu.scala 74:31]
  reg [1:0] predictor_115; // @[Bpu.scala 74:31]
  reg [1:0] predictor_116; // @[Bpu.scala 74:31]
  reg [1:0] predictor_117; // @[Bpu.scala 74:31]
  reg [1:0] predictor_118; // @[Bpu.scala 74:31]
  reg [1:0] predictor_119; // @[Bpu.scala 74:31]
  reg [1:0] predictor_120; // @[Bpu.scala 74:31]
  reg [1:0] predictor_121; // @[Bpu.scala 74:31]
  reg [1:0] predictor_122; // @[Bpu.scala 74:31]
  reg [1:0] predictor_123; // @[Bpu.scala 74:31]
  reg [1:0] predictor_124; // @[Bpu.scala 74:31]
  reg [1:0] predictor_125; // @[Bpu.scala 74:31]
  reg [1:0] predictor_126; // @[Bpu.scala 74:31]
  reg [1:0] predictor_127; // @[Bpu.scala 74:31]
  wire [31:0] _branch_mask_T = io_inst_packet_i_bits_data_0 & 32'hfc000000; // @[Lookup.scala 31:38]
  wire  _branch_mask_T_1 = 32'h10000000 == _branch_mask_T; // @[Lookup.scala 31:38]
  wire  _branch_mask_T_3 = 32'h14000000 == _branch_mask_T; // @[Lookup.scala 31:38]
  wire [31:0] _branch_mask_T_4 = io_inst_packet_i_bits_data_0 & 32'hfc1f0000; // @[Lookup.scala 31:38]
  wire  _branch_mask_T_5 = 32'h18000000 == _branch_mask_T_4; // @[Lookup.scala 31:38]
  wire  _branch_mask_T_7 = 32'h1c000000 == _branch_mask_T_4; // @[Lookup.scala 31:38]
  wire  _branch_mask_T_9 = 32'h4000000 == _branch_mask_T_4; // @[Lookup.scala 31:38]
  wire  _branch_mask_T_11 = 32'h4010000 == _branch_mask_T_4; // @[Lookup.scala 31:38]
  wire  branch_mask_0 = _branch_mask_T_1 | (_branch_mask_T_3 | (_branch_mask_T_5 | (_branch_mask_T_7 | (_branch_mask_T_9
     | (_branch_mask_T_11 | (_branch_mask_T_11 | _branch_mask_T_5)))))); // @[Lookup.scala 33:37]
  wire [31:0] _branch_mask_T_23 = io_inst_packet_i_bits_data_1 & 32'hfc000000; // @[Lookup.scala 31:38]
  wire  _branch_mask_T_24 = 32'h10000000 == _branch_mask_T_23; // @[Lookup.scala 31:38]
  wire  _branch_mask_T_26 = 32'h14000000 == _branch_mask_T_23; // @[Lookup.scala 31:38]
  wire [31:0] _branch_mask_T_27 = io_inst_packet_i_bits_data_1 & 32'hfc1f0000; // @[Lookup.scala 31:38]
  wire  _branch_mask_T_28 = 32'h18000000 == _branch_mask_T_27; // @[Lookup.scala 31:38]
  wire  _branch_mask_T_30 = 32'h1c000000 == _branch_mask_T_27; // @[Lookup.scala 31:38]
  wire  _branch_mask_T_32 = 32'h4000000 == _branch_mask_T_27; // @[Lookup.scala 31:38]
  wire  _branch_mask_T_34 = 32'h4010000 == _branch_mask_T_27; // @[Lookup.scala 31:38]
  wire  branch_mask_1 = _branch_mask_T_24 | (_branch_mask_T_26 | (_branch_mask_T_28 | (_branch_mask_T_30 | (
    _branch_mask_T_32 | (_branch_mask_T_34 | (_branch_mask_T_34 | _branch_mask_T_28)))))); // @[Lookup.scala 33:37]
  wire [31:0] _branch_mask_T_46 = io_inst_packet_i_bits_data_2 & 32'hfc000000; // @[Lookup.scala 31:38]
  wire  _branch_mask_T_47 = 32'h10000000 == _branch_mask_T_46; // @[Lookup.scala 31:38]
  wire  _branch_mask_T_49 = 32'h14000000 == _branch_mask_T_46; // @[Lookup.scala 31:38]
  wire [31:0] _branch_mask_T_50 = io_inst_packet_i_bits_data_2 & 32'hfc1f0000; // @[Lookup.scala 31:38]
  wire  _branch_mask_T_51 = 32'h18000000 == _branch_mask_T_50; // @[Lookup.scala 31:38]
  wire  _branch_mask_T_53 = 32'h1c000000 == _branch_mask_T_50; // @[Lookup.scala 31:38]
  wire  _branch_mask_T_55 = 32'h4000000 == _branch_mask_T_50; // @[Lookup.scala 31:38]
  wire  _branch_mask_T_57 = 32'h4010000 == _branch_mask_T_50; // @[Lookup.scala 31:38]
  wire  branch_mask_2 = _branch_mask_T_47 | (_branch_mask_T_49 | (_branch_mask_T_51 | (_branch_mask_T_53 | (
    _branch_mask_T_55 | (_branch_mask_T_57 | (_branch_mask_T_57 | _branch_mask_T_51)))))); // @[Lookup.scala 33:37]
  wire [31:0] _branch_mask_T_69 = io_inst_packet_i_bits_data_3 & 32'hfc000000; // @[Lookup.scala 31:38]
  wire  _branch_mask_T_70 = 32'h10000000 == _branch_mask_T_69; // @[Lookup.scala 31:38]
  wire  _branch_mask_T_72 = 32'h14000000 == _branch_mask_T_69; // @[Lookup.scala 31:38]
  wire [31:0] _branch_mask_T_73 = io_inst_packet_i_bits_data_3 & 32'hfc1f0000; // @[Lookup.scala 31:38]
  wire  _branch_mask_T_74 = 32'h18000000 == _branch_mask_T_73; // @[Lookup.scala 31:38]
  wire  _branch_mask_T_76 = 32'h1c000000 == _branch_mask_T_73; // @[Lookup.scala 31:38]
  wire  _branch_mask_T_78 = 32'h4000000 == _branch_mask_T_73; // @[Lookup.scala 31:38]
  wire  _branch_mask_T_80 = 32'h4010000 == _branch_mask_T_73; // @[Lookup.scala 31:38]
  wire  branch_mask_3 = _branch_mask_T_70 | (_branch_mask_T_72 | (_branch_mask_T_74 | (_branch_mask_T_76 | (
    _branch_mask_T_78 | (_branch_mask_T_80 | (_branch_mask_T_80 | _branch_mask_T_74)))))); // @[Lookup.scala 33:37]
  wire [31:0] _branch_mask_T_92 = io_inst_packet_i_bits_data_4 & 32'hfc000000; // @[Lookup.scala 31:38]
  wire  _branch_mask_T_93 = 32'h10000000 == _branch_mask_T_92; // @[Lookup.scala 31:38]
  wire  _branch_mask_T_95 = 32'h14000000 == _branch_mask_T_92; // @[Lookup.scala 31:38]
  wire [31:0] _branch_mask_T_96 = io_inst_packet_i_bits_data_4 & 32'hfc1f0000; // @[Lookup.scala 31:38]
  wire  _branch_mask_T_97 = 32'h18000000 == _branch_mask_T_96; // @[Lookup.scala 31:38]
  wire  _branch_mask_T_99 = 32'h1c000000 == _branch_mask_T_96; // @[Lookup.scala 31:38]
  wire  _branch_mask_T_101 = 32'h4000000 == _branch_mask_T_96; // @[Lookup.scala 31:38]
  wire  _branch_mask_T_103 = 32'h4010000 == _branch_mask_T_96; // @[Lookup.scala 31:38]
  wire  branch_mask_4 = _branch_mask_T_93 | (_branch_mask_T_95 | (_branch_mask_T_97 | (_branch_mask_T_99 | (
    _branch_mask_T_101 | (_branch_mask_T_103 | (_branch_mask_T_103 | _branch_mask_T_97)))))); // @[Lookup.scala 33:37]
  wire [31:0] _branch_mask_T_115 = io_inst_packet_i_bits_data_5 & 32'hfc000000; // @[Lookup.scala 31:38]
  wire  _branch_mask_T_116 = 32'h10000000 == _branch_mask_T_115; // @[Lookup.scala 31:38]
  wire  _branch_mask_T_118 = 32'h14000000 == _branch_mask_T_115; // @[Lookup.scala 31:38]
  wire [31:0] _branch_mask_T_119 = io_inst_packet_i_bits_data_5 & 32'hfc1f0000; // @[Lookup.scala 31:38]
  wire  _branch_mask_T_120 = 32'h18000000 == _branch_mask_T_119; // @[Lookup.scala 31:38]
  wire  _branch_mask_T_122 = 32'h1c000000 == _branch_mask_T_119; // @[Lookup.scala 31:38]
  wire  _branch_mask_T_124 = 32'h4000000 == _branch_mask_T_119; // @[Lookup.scala 31:38]
  wire  _branch_mask_T_126 = 32'h4010000 == _branch_mask_T_119; // @[Lookup.scala 31:38]
  wire  branch_mask_5 = _branch_mask_T_116 | (_branch_mask_T_118 | (_branch_mask_T_120 | (_branch_mask_T_122 | (
    _branch_mask_T_124 | (_branch_mask_T_126 | (_branch_mask_T_126 | _branch_mask_T_120)))))); // @[Lookup.scala 33:37]
  wire [31:0] _branch_mask_T_138 = io_inst_packet_i_bits_data_6 & 32'hfc000000; // @[Lookup.scala 31:38]
  wire  _branch_mask_T_139 = 32'h10000000 == _branch_mask_T_138; // @[Lookup.scala 31:38]
  wire  _branch_mask_T_141 = 32'h14000000 == _branch_mask_T_138; // @[Lookup.scala 31:38]
  wire [31:0] _branch_mask_T_142 = io_inst_packet_i_bits_data_6 & 32'hfc1f0000; // @[Lookup.scala 31:38]
  wire  _branch_mask_T_143 = 32'h18000000 == _branch_mask_T_142; // @[Lookup.scala 31:38]
  wire  _branch_mask_T_145 = 32'h1c000000 == _branch_mask_T_142; // @[Lookup.scala 31:38]
  wire  _branch_mask_T_147 = 32'h4000000 == _branch_mask_T_142; // @[Lookup.scala 31:38]
  wire  _branch_mask_T_149 = 32'h4010000 == _branch_mask_T_142; // @[Lookup.scala 31:38]
  wire  branch_mask_6 = _branch_mask_T_139 | (_branch_mask_T_141 | (_branch_mask_T_143 | (_branch_mask_T_145 | (
    _branch_mask_T_147 | (_branch_mask_T_149 | (_branch_mask_T_149 | _branch_mask_T_143)))))); // @[Lookup.scala 33:37]
  wire [31:0] _branch_mask_T_161 = io_inst_packet_i_bits_data_7 & 32'hfc000000; // @[Lookup.scala 31:38]
  wire  _branch_mask_T_162 = 32'h10000000 == _branch_mask_T_161; // @[Lookup.scala 31:38]
  wire  _branch_mask_T_164 = 32'h14000000 == _branch_mask_T_161; // @[Lookup.scala 31:38]
  wire [31:0] _branch_mask_T_165 = io_inst_packet_i_bits_data_7 & 32'hfc1f0000; // @[Lookup.scala 31:38]
  wire  _branch_mask_T_166 = 32'h18000000 == _branch_mask_T_165; // @[Lookup.scala 31:38]
  wire  _branch_mask_T_168 = 32'h1c000000 == _branch_mask_T_165; // @[Lookup.scala 31:38]
  wire  _branch_mask_T_170 = 32'h4000000 == _branch_mask_T_165; // @[Lookup.scala 31:38]
  wire  _branch_mask_T_172 = 32'h4010000 == _branch_mask_T_165; // @[Lookup.scala 31:38]
  wire  branch_mask_7 = _branch_mask_T_162 | (_branch_mask_T_164 | (_branch_mask_T_166 | (_branch_mask_T_168 | (
    _branch_mask_T_170 | (_branch_mask_T_172 | (_branch_mask_T_172 | _branch_mask_T_166)))))); // @[Lookup.scala 33:37]
  wire [7:0] _fetched_mask_T_1 = 8'h1 << io_inst_packet_i_bits_addr[4:2]; // @[OneHot.scala 58:35]
  wire  _fetched_mask_T_11 = _fetched_mask_T_1[0] | _fetched_mask_T_1[1]; // @[Bpu.scala 89:160]
  wire  _fetched_mask_T_12 = _fetched_mask_T_1[0] | _fetched_mask_T_1[1] | _fetched_mask_T_1[2]; // @[Bpu.scala 89:160]
  wire  _fetched_mask_T_13 = _fetched_mask_T_1[0] | _fetched_mask_T_1[1] | _fetched_mask_T_1[2] | _fetched_mask_T_1[3]; // @[Bpu.scala 89:160]
  wire  _fetched_mask_T_14 = _fetched_mask_T_1[0] | _fetched_mask_T_1[1] | _fetched_mask_T_1[2] | _fetched_mask_T_1[3]
     | _fetched_mask_T_1[4]; // @[Bpu.scala 89:160]
  wire  _fetched_mask_T_15 = _fetched_mask_T_1[0] | _fetched_mask_T_1[1] | _fetched_mask_T_1[2] | _fetched_mask_T_1[3]
     | _fetched_mask_T_1[4] | _fetched_mask_T_1[5]; // @[Bpu.scala 89:160]
  wire  _fetched_mask_T_16 = _fetched_mask_T_1[0] | _fetched_mask_T_1[1] | _fetched_mask_T_1[2] | _fetched_mask_T_1[3]
     | _fetched_mask_T_1[4] | _fetched_mask_T_1[5] | _fetched_mask_T_1[6]; // @[Bpu.scala 89:160]
  wire  _fetched_mask_T_17 = _fetched_mask_T_1[0] | _fetched_mask_T_1[1] | _fetched_mask_T_1[2] | _fetched_mask_T_1[3]
     | _fetched_mask_T_1[4] | _fetched_mask_T_1[5] | _fetched_mask_T_1[6] | _fetched_mask_T_1[7]; // @[Bpu.scala 89:160]
  wire [7:0] _fetched_mask_T_18 = {_fetched_mask_T_17,_fetched_mask_T_16,_fetched_mask_T_15,_fetched_mask_T_14,
    _fetched_mask_T_13,_fetched_mask_T_12,_fetched_mask_T_11,_fetched_mask_T_1[0]}; // @[Bpu.scala 89:180]
  wire [7:0] _fetched_mask_T_19 = io_is_delay ? 8'h1 : _fetched_mask_T_18; // @[Bpu.scala 89:25]
  wire  fetched_mask_0 = _fetched_mask_T_19[0]; // @[Bpu.scala 89:191]
  wire  fetched_mask_1 = _fetched_mask_T_19[1]; // @[Bpu.scala 89:191]
  wire  fetched_mask_2 = _fetched_mask_T_19[2]; // @[Bpu.scala 89:191]
  wire  fetched_mask_3 = _fetched_mask_T_19[3]; // @[Bpu.scala 89:191]
  wire  fetched_mask_4 = _fetched_mask_T_19[4]; // @[Bpu.scala 89:191]
  wire  fetched_mask_5 = _fetched_mask_T_19[5]; // @[Bpu.scala 89:191]
  wire  fetched_mask_6 = _fetched_mask_T_19[6]; // @[Bpu.scala 89:191]
  wire  fetched_mask_7 = _fetched_mask_T_19[7]; // @[Bpu.scala 89:191]
  wire  need_predict_0 = branch_mask_0 & fetched_mask_0; // @[Bpu.scala 91:67]
  wire  need_predict_1 = branch_mask_1 & fetched_mask_1; // @[Bpu.scala 91:67]
  wire  need_predict_2 = branch_mask_2 & fetched_mask_2; // @[Bpu.scala 91:67]
  wire  need_predict_3 = branch_mask_3 & fetched_mask_3; // @[Bpu.scala 91:67]
  wire  need_predict_4 = branch_mask_4 & fetched_mask_4; // @[Bpu.scala 91:67]
  wire  need_predict_5 = branch_mask_5 & fetched_mask_5; // @[Bpu.scala 91:67]
  wire  need_predict_6 = branch_mask_6 & fetched_mask_6; // @[Bpu.scala 91:67]
  wire  need_predict_7 = branch_mask_7 & fetched_mask_7; // @[Bpu.scala 91:67]
  wire  predictor_idx_hi_lo = io_inst_packet_i_bits_addr[5]; // @[Bpu.scala 94:66]
  wire [7:0] predictor_idx_0 = {global_history,predictor_idx_hi_lo,3'h0}; // @[Cat.scala 30:58]
  wire [7:0] predictor_idx_1 = {global_history,predictor_idx_hi_lo,3'h1}; // @[Cat.scala 30:58]
  wire [7:0] predictor_idx_2 = {global_history,predictor_idx_hi_lo,3'h2}; // @[Cat.scala 30:58]
  wire [7:0] predictor_idx_3 = {global_history,predictor_idx_hi_lo,3'h3}; // @[Cat.scala 30:58]
  wire [7:0] predictor_idx_4 = {global_history,predictor_idx_hi_lo,3'h4}; // @[Cat.scala 30:58]
  wire [7:0] predictor_idx_5 = {global_history,predictor_idx_hi_lo,3'h5}; // @[Cat.scala 30:58]
  wire [7:0] predictor_idx_6 = {global_history,predictor_idx_hi_lo,3'h6}; // @[Cat.scala 30:58]
  wire [7:0] predictor_idx_7 = {global_history,predictor_idx_hi_lo,3'h7}; // @[Cat.scala 30:58]
  wire [1:0] _GEN_1 = 7'h1 == predictor_idx_0[6:0] ? predictor_1 : predictor_0; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_2 = 7'h2 == predictor_idx_0[6:0] ? predictor_2 : _GEN_1; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_3 = 7'h3 == predictor_idx_0[6:0] ? predictor_3 : _GEN_2; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_4 = 7'h4 == predictor_idx_0[6:0] ? predictor_4 : _GEN_3; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_5 = 7'h5 == predictor_idx_0[6:0] ? predictor_5 : _GEN_4; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_6 = 7'h6 == predictor_idx_0[6:0] ? predictor_6 : _GEN_5; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_7 = 7'h7 == predictor_idx_0[6:0] ? predictor_7 : _GEN_6; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_8 = 7'h8 == predictor_idx_0[6:0] ? predictor_8 : _GEN_7; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_9 = 7'h9 == predictor_idx_0[6:0] ? predictor_9 : _GEN_8; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_10 = 7'ha == predictor_idx_0[6:0] ? predictor_10 : _GEN_9; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_11 = 7'hb == predictor_idx_0[6:0] ? predictor_11 : _GEN_10; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_12 = 7'hc == predictor_idx_0[6:0] ? predictor_12 : _GEN_11; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_13 = 7'hd == predictor_idx_0[6:0] ? predictor_13 : _GEN_12; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_14 = 7'he == predictor_idx_0[6:0] ? predictor_14 : _GEN_13; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_15 = 7'hf == predictor_idx_0[6:0] ? predictor_15 : _GEN_14; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_16 = 7'h10 == predictor_idx_0[6:0] ? predictor_16 : _GEN_15; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_17 = 7'h11 == predictor_idx_0[6:0] ? predictor_17 : _GEN_16; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_18 = 7'h12 == predictor_idx_0[6:0] ? predictor_18 : _GEN_17; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_19 = 7'h13 == predictor_idx_0[6:0] ? predictor_19 : _GEN_18; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_20 = 7'h14 == predictor_idx_0[6:0] ? predictor_20 : _GEN_19; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_21 = 7'h15 == predictor_idx_0[6:0] ? predictor_21 : _GEN_20; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_22 = 7'h16 == predictor_idx_0[6:0] ? predictor_22 : _GEN_21; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_23 = 7'h17 == predictor_idx_0[6:0] ? predictor_23 : _GEN_22; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_24 = 7'h18 == predictor_idx_0[6:0] ? predictor_24 : _GEN_23; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_25 = 7'h19 == predictor_idx_0[6:0] ? predictor_25 : _GEN_24; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_26 = 7'h1a == predictor_idx_0[6:0] ? predictor_26 : _GEN_25; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_27 = 7'h1b == predictor_idx_0[6:0] ? predictor_27 : _GEN_26; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_28 = 7'h1c == predictor_idx_0[6:0] ? predictor_28 : _GEN_27; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_29 = 7'h1d == predictor_idx_0[6:0] ? predictor_29 : _GEN_28; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_30 = 7'h1e == predictor_idx_0[6:0] ? predictor_30 : _GEN_29; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_31 = 7'h1f == predictor_idx_0[6:0] ? predictor_31 : _GEN_30; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_32 = 7'h20 == predictor_idx_0[6:0] ? predictor_32 : _GEN_31; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_33 = 7'h21 == predictor_idx_0[6:0] ? predictor_33 : _GEN_32; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_34 = 7'h22 == predictor_idx_0[6:0] ? predictor_34 : _GEN_33; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_35 = 7'h23 == predictor_idx_0[6:0] ? predictor_35 : _GEN_34; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_36 = 7'h24 == predictor_idx_0[6:0] ? predictor_36 : _GEN_35; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_37 = 7'h25 == predictor_idx_0[6:0] ? predictor_37 : _GEN_36; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_38 = 7'h26 == predictor_idx_0[6:0] ? predictor_38 : _GEN_37; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_39 = 7'h27 == predictor_idx_0[6:0] ? predictor_39 : _GEN_38; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_40 = 7'h28 == predictor_idx_0[6:0] ? predictor_40 : _GEN_39; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_41 = 7'h29 == predictor_idx_0[6:0] ? predictor_41 : _GEN_40; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_42 = 7'h2a == predictor_idx_0[6:0] ? predictor_42 : _GEN_41; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_43 = 7'h2b == predictor_idx_0[6:0] ? predictor_43 : _GEN_42; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_44 = 7'h2c == predictor_idx_0[6:0] ? predictor_44 : _GEN_43; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_45 = 7'h2d == predictor_idx_0[6:0] ? predictor_45 : _GEN_44; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_46 = 7'h2e == predictor_idx_0[6:0] ? predictor_46 : _GEN_45; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_47 = 7'h2f == predictor_idx_0[6:0] ? predictor_47 : _GEN_46; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_48 = 7'h30 == predictor_idx_0[6:0] ? predictor_48 : _GEN_47; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_49 = 7'h31 == predictor_idx_0[6:0] ? predictor_49 : _GEN_48; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_50 = 7'h32 == predictor_idx_0[6:0] ? predictor_50 : _GEN_49; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_51 = 7'h33 == predictor_idx_0[6:0] ? predictor_51 : _GEN_50; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_52 = 7'h34 == predictor_idx_0[6:0] ? predictor_52 : _GEN_51; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_53 = 7'h35 == predictor_idx_0[6:0] ? predictor_53 : _GEN_52; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_54 = 7'h36 == predictor_idx_0[6:0] ? predictor_54 : _GEN_53; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_55 = 7'h37 == predictor_idx_0[6:0] ? predictor_55 : _GEN_54; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_56 = 7'h38 == predictor_idx_0[6:0] ? predictor_56 : _GEN_55; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_57 = 7'h39 == predictor_idx_0[6:0] ? predictor_57 : _GEN_56; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_58 = 7'h3a == predictor_idx_0[6:0] ? predictor_58 : _GEN_57; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_59 = 7'h3b == predictor_idx_0[6:0] ? predictor_59 : _GEN_58; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_60 = 7'h3c == predictor_idx_0[6:0] ? predictor_60 : _GEN_59; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_61 = 7'h3d == predictor_idx_0[6:0] ? predictor_61 : _GEN_60; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_62 = 7'h3e == predictor_idx_0[6:0] ? predictor_62 : _GEN_61; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_63 = 7'h3f == predictor_idx_0[6:0] ? predictor_63 : _GEN_62; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_64 = 7'h40 == predictor_idx_0[6:0] ? predictor_64 : _GEN_63; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_65 = 7'h41 == predictor_idx_0[6:0] ? predictor_65 : _GEN_64; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_66 = 7'h42 == predictor_idx_0[6:0] ? predictor_66 : _GEN_65; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_67 = 7'h43 == predictor_idx_0[6:0] ? predictor_67 : _GEN_66; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_68 = 7'h44 == predictor_idx_0[6:0] ? predictor_68 : _GEN_67; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_69 = 7'h45 == predictor_idx_0[6:0] ? predictor_69 : _GEN_68; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_70 = 7'h46 == predictor_idx_0[6:0] ? predictor_70 : _GEN_69; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_71 = 7'h47 == predictor_idx_0[6:0] ? predictor_71 : _GEN_70; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_72 = 7'h48 == predictor_idx_0[6:0] ? predictor_72 : _GEN_71; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_73 = 7'h49 == predictor_idx_0[6:0] ? predictor_73 : _GEN_72; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_74 = 7'h4a == predictor_idx_0[6:0] ? predictor_74 : _GEN_73; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_75 = 7'h4b == predictor_idx_0[6:0] ? predictor_75 : _GEN_74; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_76 = 7'h4c == predictor_idx_0[6:0] ? predictor_76 : _GEN_75; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_77 = 7'h4d == predictor_idx_0[6:0] ? predictor_77 : _GEN_76; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_78 = 7'h4e == predictor_idx_0[6:0] ? predictor_78 : _GEN_77; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_79 = 7'h4f == predictor_idx_0[6:0] ? predictor_79 : _GEN_78; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_80 = 7'h50 == predictor_idx_0[6:0] ? predictor_80 : _GEN_79; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_81 = 7'h51 == predictor_idx_0[6:0] ? predictor_81 : _GEN_80; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_82 = 7'h52 == predictor_idx_0[6:0] ? predictor_82 : _GEN_81; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_83 = 7'h53 == predictor_idx_0[6:0] ? predictor_83 : _GEN_82; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_84 = 7'h54 == predictor_idx_0[6:0] ? predictor_84 : _GEN_83; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_85 = 7'h55 == predictor_idx_0[6:0] ? predictor_85 : _GEN_84; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_86 = 7'h56 == predictor_idx_0[6:0] ? predictor_86 : _GEN_85; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_87 = 7'h57 == predictor_idx_0[6:0] ? predictor_87 : _GEN_86; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_88 = 7'h58 == predictor_idx_0[6:0] ? predictor_88 : _GEN_87; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_89 = 7'h59 == predictor_idx_0[6:0] ? predictor_89 : _GEN_88; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_90 = 7'h5a == predictor_idx_0[6:0] ? predictor_90 : _GEN_89; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_91 = 7'h5b == predictor_idx_0[6:0] ? predictor_91 : _GEN_90; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_92 = 7'h5c == predictor_idx_0[6:0] ? predictor_92 : _GEN_91; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_93 = 7'h5d == predictor_idx_0[6:0] ? predictor_93 : _GEN_92; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_94 = 7'h5e == predictor_idx_0[6:0] ? predictor_94 : _GEN_93; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_95 = 7'h5f == predictor_idx_0[6:0] ? predictor_95 : _GEN_94; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_96 = 7'h60 == predictor_idx_0[6:0] ? predictor_96 : _GEN_95; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_97 = 7'h61 == predictor_idx_0[6:0] ? predictor_97 : _GEN_96; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_98 = 7'h62 == predictor_idx_0[6:0] ? predictor_98 : _GEN_97; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_99 = 7'h63 == predictor_idx_0[6:0] ? predictor_99 : _GEN_98; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_100 = 7'h64 == predictor_idx_0[6:0] ? predictor_100 : _GEN_99; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_101 = 7'h65 == predictor_idx_0[6:0] ? predictor_101 : _GEN_100; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_102 = 7'h66 == predictor_idx_0[6:0] ? predictor_102 : _GEN_101; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_103 = 7'h67 == predictor_idx_0[6:0] ? predictor_103 : _GEN_102; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_104 = 7'h68 == predictor_idx_0[6:0] ? predictor_104 : _GEN_103; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_105 = 7'h69 == predictor_idx_0[6:0] ? predictor_105 : _GEN_104; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_106 = 7'h6a == predictor_idx_0[6:0] ? predictor_106 : _GEN_105; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_107 = 7'h6b == predictor_idx_0[6:0] ? predictor_107 : _GEN_106; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_108 = 7'h6c == predictor_idx_0[6:0] ? predictor_108 : _GEN_107; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_109 = 7'h6d == predictor_idx_0[6:0] ? predictor_109 : _GEN_108; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_110 = 7'h6e == predictor_idx_0[6:0] ? predictor_110 : _GEN_109; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_111 = 7'h6f == predictor_idx_0[6:0] ? predictor_111 : _GEN_110; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_112 = 7'h70 == predictor_idx_0[6:0] ? predictor_112 : _GEN_111; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_113 = 7'h71 == predictor_idx_0[6:0] ? predictor_113 : _GEN_112; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_114 = 7'h72 == predictor_idx_0[6:0] ? predictor_114 : _GEN_113; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_115 = 7'h73 == predictor_idx_0[6:0] ? predictor_115 : _GEN_114; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_116 = 7'h74 == predictor_idx_0[6:0] ? predictor_116 : _GEN_115; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_117 = 7'h75 == predictor_idx_0[6:0] ? predictor_117 : _GEN_116; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_118 = 7'h76 == predictor_idx_0[6:0] ? predictor_118 : _GEN_117; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_119 = 7'h77 == predictor_idx_0[6:0] ? predictor_119 : _GEN_118; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_120 = 7'h78 == predictor_idx_0[6:0] ? predictor_120 : _GEN_119; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_121 = 7'h79 == predictor_idx_0[6:0] ? predictor_121 : _GEN_120; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_122 = 7'h7a == predictor_idx_0[6:0] ? predictor_122 : _GEN_121; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_123 = 7'h7b == predictor_idx_0[6:0] ? predictor_123 : _GEN_122; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_124 = 7'h7c == predictor_idx_0[6:0] ? predictor_124 : _GEN_123; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_125 = 7'h7d == predictor_idx_0[6:0] ? predictor_125 : _GEN_124; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_126 = 7'h7e == predictor_idx_0[6:0] ? predictor_126 : _GEN_125; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_127 = 7'h7f == predictor_idx_0[6:0] ? predictor_127 : _GEN_126; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire  predict_mask_0 = _GEN_127[1]; // @[Bpu.scala 96:62]
  wire [1:0] _GEN_129 = 7'h1 == predictor_idx_1[6:0] ? predictor_1 : predictor_0; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_130 = 7'h2 == predictor_idx_1[6:0] ? predictor_2 : _GEN_129; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_131 = 7'h3 == predictor_idx_1[6:0] ? predictor_3 : _GEN_130; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_132 = 7'h4 == predictor_idx_1[6:0] ? predictor_4 : _GEN_131; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_133 = 7'h5 == predictor_idx_1[6:0] ? predictor_5 : _GEN_132; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_134 = 7'h6 == predictor_idx_1[6:0] ? predictor_6 : _GEN_133; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_135 = 7'h7 == predictor_idx_1[6:0] ? predictor_7 : _GEN_134; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_136 = 7'h8 == predictor_idx_1[6:0] ? predictor_8 : _GEN_135; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_137 = 7'h9 == predictor_idx_1[6:0] ? predictor_9 : _GEN_136; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_138 = 7'ha == predictor_idx_1[6:0] ? predictor_10 : _GEN_137; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_139 = 7'hb == predictor_idx_1[6:0] ? predictor_11 : _GEN_138; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_140 = 7'hc == predictor_idx_1[6:0] ? predictor_12 : _GEN_139; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_141 = 7'hd == predictor_idx_1[6:0] ? predictor_13 : _GEN_140; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_142 = 7'he == predictor_idx_1[6:0] ? predictor_14 : _GEN_141; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_143 = 7'hf == predictor_idx_1[6:0] ? predictor_15 : _GEN_142; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_144 = 7'h10 == predictor_idx_1[6:0] ? predictor_16 : _GEN_143; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_145 = 7'h11 == predictor_idx_1[6:0] ? predictor_17 : _GEN_144; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_146 = 7'h12 == predictor_idx_1[6:0] ? predictor_18 : _GEN_145; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_147 = 7'h13 == predictor_idx_1[6:0] ? predictor_19 : _GEN_146; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_148 = 7'h14 == predictor_idx_1[6:0] ? predictor_20 : _GEN_147; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_149 = 7'h15 == predictor_idx_1[6:0] ? predictor_21 : _GEN_148; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_150 = 7'h16 == predictor_idx_1[6:0] ? predictor_22 : _GEN_149; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_151 = 7'h17 == predictor_idx_1[6:0] ? predictor_23 : _GEN_150; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_152 = 7'h18 == predictor_idx_1[6:0] ? predictor_24 : _GEN_151; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_153 = 7'h19 == predictor_idx_1[6:0] ? predictor_25 : _GEN_152; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_154 = 7'h1a == predictor_idx_1[6:0] ? predictor_26 : _GEN_153; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_155 = 7'h1b == predictor_idx_1[6:0] ? predictor_27 : _GEN_154; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_156 = 7'h1c == predictor_idx_1[6:0] ? predictor_28 : _GEN_155; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_157 = 7'h1d == predictor_idx_1[6:0] ? predictor_29 : _GEN_156; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_158 = 7'h1e == predictor_idx_1[6:0] ? predictor_30 : _GEN_157; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_159 = 7'h1f == predictor_idx_1[6:0] ? predictor_31 : _GEN_158; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_160 = 7'h20 == predictor_idx_1[6:0] ? predictor_32 : _GEN_159; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_161 = 7'h21 == predictor_idx_1[6:0] ? predictor_33 : _GEN_160; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_162 = 7'h22 == predictor_idx_1[6:0] ? predictor_34 : _GEN_161; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_163 = 7'h23 == predictor_idx_1[6:0] ? predictor_35 : _GEN_162; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_164 = 7'h24 == predictor_idx_1[6:0] ? predictor_36 : _GEN_163; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_165 = 7'h25 == predictor_idx_1[6:0] ? predictor_37 : _GEN_164; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_166 = 7'h26 == predictor_idx_1[6:0] ? predictor_38 : _GEN_165; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_167 = 7'h27 == predictor_idx_1[6:0] ? predictor_39 : _GEN_166; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_168 = 7'h28 == predictor_idx_1[6:0] ? predictor_40 : _GEN_167; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_169 = 7'h29 == predictor_idx_1[6:0] ? predictor_41 : _GEN_168; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_170 = 7'h2a == predictor_idx_1[6:0] ? predictor_42 : _GEN_169; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_171 = 7'h2b == predictor_idx_1[6:0] ? predictor_43 : _GEN_170; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_172 = 7'h2c == predictor_idx_1[6:0] ? predictor_44 : _GEN_171; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_173 = 7'h2d == predictor_idx_1[6:0] ? predictor_45 : _GEN_172; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_174 = 7'h2e == predictor_idx_1[6:0] ? predictor_46 : _GEN_173; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_175 = 7'h2f == predictor_idx_1[6:0] ? predictor_47 : _GEN_174; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_176 = 7'h30 == predictor_idx_1[6:0] ? predictor_48 : _GEN_175; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_177 = 7'h31 == predictor_idx_1[6:0] ? predictor_49 : _GEN_176; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_178 = 7'h32 == predictor_idx_1[6:0] ? predictor_50 : _GEN_177; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_179 = 7'h33 == predictor_idx_1[6:0] ? predictor_51 : _GEN_178; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_180 = 7'h34 == predictor_idx_1[6:0] ? predictor_52 : _GEN_179; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_181 = 7'h35 == predictor_idx_1[6:0] ? predictor_53 : _GEN_180; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_182 = 7'h36 == predictor_idx_1[6:0] ? predictor_54 : _GEN_181; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_183 = 7'h37 == predictor_idx_1[6:0] ? predictor_55 : _GEN_182; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_184 = 7'h38 == predictor_idx_1[6:0] ? predictor_56 : _GEN_183; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_185 = 7'h39 == predictor_idx_1[6:0] ? predictor_57 : _GEN_184; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_186 = 7'h3a == predictor_idx_1[6:0] ? predictor_58 : _GEN_185; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_187 = 7'h3b == predictor_idx_1[6:0] ? predictor_59 : _GEN_186; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_188 = 7'h3c == predictor_idx_1[6:0] ? predictor_60 : _GEN_187; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_189 = 7'h3d == predictor_idx_1[6:0] ? predictor_61 : _GEN_188; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_190 = 7'h3e == predictor_idx_1[6:0] ? predictor_62 : _GEN_189; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_191 = 7'h3f == predictor_idx_1[6:0] ? predictor_63 : _GEN_190; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_192 = 7'h40 == predictor_idx_1[6:0] ? predictor_64 : _GEN_191; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_193 = 7'h41 == predictor_idx_1[6:0] ? predictor_65 : _GEN_192; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_194 = 7'h42 == predictor_idx_1[6:0] ? predictor_66 : _GEN_193; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_195 = 7'h43 == predictor_idx_1[6:0] ? predictor_67 : _GEN_194; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_196 = 7'h44 == predictor_idx_1[6:0] ? predictor_68 : _GEN_195; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_197 = 7'h45 == predictor_idx_1[6:0] ? predictor_69 : _GEN_196; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_198 = 7'h46 == predictor_idx_1[6:0] ? predictor_70 : _GEN_197; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_199 = 7'h47 == predictor_idx_1[6:0] ? predictor_71 : _GEN_198; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_200 = 7'h48 == predictor_idx_1[6:0] ? predictor_72 : _GEN_199; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_201 = 7'h49 == predictor_idx_1[6:0] ? predictor_73 : _GEN_200; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_202 = 7'h4a == predictor_idx_1[6:0] ? predictor_74 : _GEN_201; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_203 = 7'h4b == predictor_idx_1[6:0] ? predictor_75 : _GEN_202; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_204 = 7'h4c == predictor_idx_1[6:0] ? predictor_76 : _GEN_203; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_205 = 7'h4d == predictor_idx_1[6:0] ? predictor_77 : _GEN_204; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_206 = 7'h4e == predictor_idx_1[6:0] ? predictor_78 : _GEN_205; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_207 = 7'h4f == predictor_idx_1[6:0] ? predictor_79 : _GEN_206; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_208 = 7'h50 == predictor_idx_1[6:0] ? predictor_80 : _GEN_207; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_209 = 7'h51 == predictor_idx_1[6:0] ? predictor_81 : _GEN_208; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_210 = 7'h52 == predictor_idx_1[6:0] ? predictor_82 : _GEN_209; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_211 = 7'h53 == predictor_idx_1[6:0] ? predictor_83 : _GEN_210; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_212 = 7'h54 == predictor_idx_1[6:0] ? predictor_84 : _GEN_211; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_213 = 7'h55 == predictor_idx_1[6:0] ? predictor_85 : _GEN_212; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_214 = 7'h56 == predictor_idx_1[6:0] ? predictor_86 : _GEN_213; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_215 = 7'h57 == predictor_idx_1[6:0] ? predictor_87 : _GEN_214; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_216 = 7'h58 == predictor_idx_1[6:0] ? predictor_88 : _GEN_215; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_217 = 7'h59 == predictor_idx_1[6:0] ? predictor_89 : _GEN_216; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_218 = 7'h5a == predictor_idx_1[6:0] ? predictor_90 : _GEN_217; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_219 = 7'h5b == predictor_idx_1[6:0] ? predictor_91 : _GEN_218; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_220 = 7'h5c == predictor_idx_1[6:0] ? predictor_92 : _GEN_219; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_221 = 7'h5d == predictor_idx_1[6:0] ? predictor_93 : _GEN_220; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_222 = 7'h5e == predictor_idx_1[6:0] ? predictor_94 : _GEN_221; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_223 = 7'h5f == predictor_idx_1[6:0] ? predictor_95 : _GEN_222; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_224 = 7'h60 == predictor_idx_1[6:0] ? predictor_96 : _GEN_223; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_225 = 7'h61 == predictor_idx_1[6:0] ? predictor_97 : _GEN_224; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_226 = 7'h62 == predictor_idx_1[6:0] ? predictor_98 : _GEN_225; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_227 = 7'h63 == predictor_idx_1[6:0] ? predictor_99 : _GEN_226; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_228 = 7'h64 == predictor_idx_1[6:0] ? predictor_100 : _GEN_227; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_229 = 7'h65 == predictor_idx_1[6:0] ? predictor_101 : _GEN_228; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_230 = 7'h66 == predictor_idx_1[6:0] ? predictor_102 : _GEN_229; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_231 = 7'h67 == predictor_idx_1[6:0] ? predictor_103 : _GEN_230; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_232 = 7'h68 == predictor_idx_1[6:0] ? predictor_104 : _GEN_231; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_233 = 7'h69 == predictor_idx_1[6:0] ? predictor_105 : _GEN_232; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_234 = 7'h6a == predictor_idx_1[6:0] ? predictor_106 : _GEN_233; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_235 = 7'h6b == predictor_idx_1[6:0] ? predictor_107 : _GEN_234; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_236 = 7'h6c == predictor_idx_1[6:0] ? predictor_108 : _GEN_235; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_237 = 7'h6d == predictor_idx_1[6:0] ? predictor_109 : _GEN_236; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_238 = 7'h6e == predictor_idx_1[6:0] ? predictor_110 : _GEN_237; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_239 = 7'h6f == predictor_idx_1[6:0] ? predictor_111 : _GEN_238; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_240 = 7'h70 == predictor_idx_1[6:0] ? predictor_112 : _GEN_239; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_241 = 7'h71 == predictor_idx_1[6:0] ? predictor_113 : _GEN_240; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_242 = 7'h72 == predictor_idx_1[6:0] ? predictor_114 : _GEN_241; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_243 = 7'h73 == predictor_idx_1[6:0] ? predictor_115 : _GEN_242; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_244 = 7'h74 == predictor_idx_1[6:0] ? predictor_116 : _GEN_243; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_245 = 7'h75 == predictor_idx_1[6:0] ? predictor_117 : _GEN_244; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_246 = 7'h76 == predictor_idx_1[6:0] ? predictor_118 : _GEN_245; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_247 = 7'h77 == predictor_idx_1[6:0] ? predictor_119 : _GEN_246; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_248 = 7'h78 == predictor_idx_1[6:0] ? predictor_120 : _GEN_247; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_249 = 7'h79 == predictor_idx_1[6:0] ? predictor_121 : _GEN_248; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_250 = 7'h7a == predictor_idx_1[6:0] ? predictor_122 : _GEN_249; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_251 = 7'h7b == predictor_idx_1[6:0] ? predictor_123 : _GEN_250; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_252 = 7'h7c == predictor_idx_1[6:0] ? predictor_124 : _GEN_251; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_253 = 7'h7d == predictor_idx_1[6:0] ? predictor_125 : _GEN_252; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_254 = 7'h7e == predictor_idx_1[6:0] ? predictor_126 : _GEN_253; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_255 = 7'h7f == predictor_idx_1[6:0] ? predictor_127 : _GEN_254; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire  predict_mask_1 = _GEN_255[1]; // @[Bpu.scala 96:62]
  wire [1:0] _GEN_257 = 7'h1 == predictor_idx_2[6:0] ? predictor_1 : predictor_0; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_258 = 7'h2 == predictor_idx_2[6:0] ? predictor_2 : _GEN_257; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_259 = 7'h3 == predictor_idx_2[6:0] ? predictor_3 : _GEN_258; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_260 = 7'h4 == predictor_idx_2[6:0] ? predictor_4 : _GEN_259; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_261 = 7'h5 == predictor_idx_2[6:0] ? predictor_5 : _GEN_260; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_262 = 7'h6 == predictor_idx_2[6:0] ? predictor_6 : _GEN_261; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_263 = 7'h7 == predictor_idx_2[6:0] ? predictor_7 : _GEN_262; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_264 = 7'h8 == predictor_idx_2[6:0] ? predictor_8 : _GEN_263; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_265 = 7'h9 == predictor_idx_2[6:0] ? predictor_9 : _GEN_264; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_266 = 7'ha == predictor_idx_2[6:0] ? predictor_10 : _GEN_265; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_267 = 7'hb == predictor_idx_2[6:0] ? predictor_11 : _GEN_266; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_268 = 7'hc == predictor_idx_2[6:0] ? predictor_12 : _GEN_267; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_269 = 7'hd == predictor_idx_2[6:0] ? predictor_13 : _GEN_268; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_270 = 7'he == predictor_idx_2[6:0] ? predictor_14 : _GEN_269; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_271 = 7'hf == predictor_idx_2[6:0] ? predictor_15 : _GEN_270; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_272 = 7'h10 == predictor_idx_2[6:0] ? predictor_16 : _GEN_271; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_273 = 7'h11 == predictor_idx_2[6:0] ? predictor_17 : _GEN_272; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_274 = 7'h12 == predictor_idx_2[6:0] ? predictor_18 : _GEN_273; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_275 = 7'h13 == predictor_idx_2[6:0] ? predictor_19 : _GEN_274; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_276 = 7'h14 == predictor_idx_2[6:0] ? predictor_20 : _GEN_275; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_277 = 7'h15 == predictor_idx_2[6:0] ? predictor_21 : _GEN_276; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_278 = 7'h16 == predictor_idx_2[6:0] ? predictor_22 : _GEN_277; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_279 = 7'h17 == predictor_idx_2[6:0] ? predictor_23 : _GEN_278; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_280 = 7'h18 == predictor_idx_2[6:0] ? predictor_24 : _GEN_279; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_281 = 7'h19 == predictor_idx_2[6:0] ? predictor_25 : _GEN_280; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_282 = 7'h1a == predictor_idx_2[6:0] ? predictor_26 : _GEN_281; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_283 = 7'h1b == predictor_idx_2[6:0] ? predictor_27 : _GEN_282; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_284 = 7'h1c == predictor_idx_2[6:0] ? predictor_28 : _GEN_283; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_285 = 7'h1d == predictor_idx_2[6:0] ? predictor_29 : _GEN_284; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_286 = 7'h1e == predictor_idx_2[6:0] ? predictor_30 : _GEN_285; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_287 = 7'h1f == predictor_idx_2[6:0] ? predictor_31 : _GEN_286; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_288 = 7'h20 == predictor_idx_2[6:0] ? predictor_32 : _GEN_287; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_289 = 7'h21 == predictor_idx_2[6:0] ? predictor_33 : _GEN_288; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_290 = 7'h22 == predictor_idx_2[6:0] ? predictor_34 : _GEN_289; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_291 = 7'h23 == predictor_idx_2[6:0] ? predictor_35 : _GEN_290; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_292 = 7'h24 == predictor_idx_2[6:0] ? predictor_36 : _GEN_291; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_293 = 7'h25 == predictor_idx_2[6:0] ? predictor_37 : _GEN_292; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_294 = 7'h26 == predictor_idx_2[6:0] ? predictor_38 : _GEN_293; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_295 = 7'h27 == predictor_idx_2[6:0] ? predictor_39 : _GEN_294; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_296 = 7'h28 == predictor_idx_2[6:0] ? predictor_40 : _GEN_295; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_297 = 7'h29 == predictor_idx_2[6:0] ? predictor_41 : _GEN_296; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_298 = 7'h2a == predictor_idx_2[6:0] ? predictor_42 : _GEN_297; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_299 = 7'h2b == predictor_idx_2[6:0] ? predictor_43 : _GEN_298; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_300 = 7'h2c == predictor_idx_2[6:0] ? predictor_44 : _GEN_299; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_301 = 7'h2d == predictor_idx_2[6:0] ? predictor_45 : _GEN_300; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_302 = 7'h2e == predictor_idx_2[6:0] ? predictor_46 : _GEN_301; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_303 = 7'h2f == predictor_idx_2[6:0] ? predictor_47 : _GEN_302; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_304 = 7'h30 == predictor_idx_2[6:0] ? predictor_48 : _GEN_303; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_305 = 7'h31 == predictor_idx_2[6:0] ? predictor_49 : _GEN_304; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_306 = 7'h32 == predictor_idx_2[6:0] ? predictor_50 : _GEN_305; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_307 = 7'h33 == predictor_idx_2[6:0] ? predictor_51 : _GEN_306; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_308 = 7'h34 == predictor_idx_2[6:0] ? predictor_52 : _GEN_307; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_309 = 7'h35 == predictor_idx_2[6:0] ? predictor_53 : _GEN_308; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_310 = 7'h36 == predictor_idx_2[6:0] ? predictor_54 : _GEN_309; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_311 = 7'h37 == predictor_idx_2[6:0] ? predictor_55 : _GEN_310; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_312 = 7'h38 == predictor_idx_2[6:0] ? predictor_56 : _GEN_311; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_313 = 7'h39 == predictor_idx_2[6:0] ? predictor_57 : _GEN_312; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_314 = 7'h3a == predictor_idx_2[6:0] ? predictor_58 : _GEN_313; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_315 = 7'h3b == predictor_idx_2[6:0] ? predictor_59 : _GEN_314; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_316 = 7'h3c == predictor_idx_2[6:0] ? predictor_60 : _GEN_315; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_317 = 7'h3d == predictor_idx_2[6:0] ? predictor_61 : _GEN_316; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_318 = 7'h3e == predictor_idx_2[6:0] ? predictor_62 : _GEN_317; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_319 = 7'h3f == predictor_idx_2[6:0] ? predictor_63 : _GEN_318; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_320 = 7'h40 == predictor_idx_2[6:0] ? predictor_64 : _GEN_319; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_321 = 7'h41 == predictor_idx_2[6:0] ? predictor_65 : _GEN_320; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_322 = 7'h42 == predictor_idx_2[6:0] ? predictor_66 : _GEN_321; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_323 = 7'h43 == predictor_idx_2[6:0] ? predictor_67 : _GEN_322; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_324 = 7'h44 == predictor_idx_2[6:0] ? predictor_68 : _GEN_323; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_325 = 7'h45 == predictor_idx_2[6:0] ? predictor_69 : _GEN_324; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_326 = 7'h46 == predictor_idx_2[6:0] ? predictor_70 : _GEN_325; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_327 = 7'h47 == predictor_idx_2[6:0] ? predictor_71 : _GEN_326; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_328 = 7'h48 == predictor_idx_2[6:0] ? predictor_72 : _GEN_327; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_329 = 7'h49 == predictor_idx_2[6:0] ? predictor_73 : _GEN_328; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_330 = 7'h4a == predictor_idx_2[6:0] ? predictor_74 : _GEN_329; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_331 = 7'h4b == predictor_idx_2[6:0] ? predictor_75 : _GEN_330; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_332 = 7'h4c == predictor_idx_2[6:0] ? predictor_76 : _GEN_331; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_333 = 7'h4d == predictor_idx_2[6:0] ? predictor_77 : _GEN_332; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_334 = 7'h4e == predictor_idx_2[6:0] ? predictor_78 : _GEN_333; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_335 = 7'h4f == predictor_idx_2[6:0] ? predictor_79 : _GEN_334; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_336 = 7'h50 == predictor_idx_2[6:0] ? predictor_80 : _GEN_335; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_337 = 7'h51 == predictor_idx_2[6:0] ? predictor_81 : _GEN_336; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_338 = 7'h52 == predictor_idx_2[6:0] ? predictor_82 : _GEN_337; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_339 = 7'h53 == predictor_idx_2[6:0] ? predictor_83 : _GEN_338; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_340 = 7'h54 == predictor_idx_2[6:0] ? predictor_84 : _GEN_339; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_341 = 7'h55 == predictor_idx_2[6:0] ? predictor_85 : _GEN_340; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_342 = 7'h56 == predictor_idx_2[6:0] ? predictor_86 : _GEN_341; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_343 = 7'h57 == predictor_idx_2[6:0] ? predictor_87 : _GEN_342; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_344 = 7'h58 == predictor_idx_2[6:0] ? predictor_88 : _GEN_343; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_345 = 7'h59 == predictor_idx_2[6:0] ? predictor_89 : _GEN_344; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_346 = 7'h5a == predictor_idx_2[6:0] ? predictor_90 : _GEN_345; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_347 = 7'h5b == predictor_idx_2[6:0] ? predictor_91 : _GEN_346; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_348 = 7'h5c == predictor_idx_2[6:0] ? predictor_92 : _GEN_347; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_349 = 7'h5d == predictor_idx_2[6:0] ? predictor_93 : _GEN_348; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_350 = 7'h5e == predictor_idx_2[6:0] ? predictor_94 : _GEN_349; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_351 = 7'h5f == predictor_idx_2[6:0] ? predictor_95 : _GEN_350; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_352 = 7'h60 == predictor_idx_2[6:0] ? predictor_96 : _GEN_351; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_353 = 7'h61 == predictor_idx_2[6:0] ? predictor_97 : _GEN_352; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_354 = 7'h62 == predictor_idx_2[6:0] ? predictor_98 : _GEN_353; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_355 = 7'h63 == predictor_idx_2[6:0] ? predictor_99 : _GEN_354; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_356 = 7'h64 == predictor_idx_2[6:0] ? predictor_100 : _GEN_355; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_357 = 7'h65 == predictor_idx_2[6:0] ? predictor_101 : _GEN_356; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_358 = 7'h66 == predictor_idx_2[6:0] ? predictor_102 : _GEN_357; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_359 = 7'h67 == predictor_idx_2[6:0] ? predictor_103 : _GEN_358; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_360 = 7'h68 == predictor_idx_2[6:0] ? predictor_104 : _GEN_359; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_361 = 7'h69 == predictor_idx_2[6:0] ? predictor_105 : _GEN_360; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_362 = 7'h6a == predictor_idx_2[6:0] ? predictor_106 : _GEN_361; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_363 = 7'h6b == predictor_idx_2[6:0] ? predictor_107 : _GEN_362; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_364 = 7'h6c == predictor_idx_2[6:0] ? predictor_108 : _GEN_363; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_365 = 7'h6d == predictor_idx_2[6:0] ? predictor_109 : _GEN_364; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_366 = 7'h6e == predictor_idx_2[6:0] ? predictor_110 : _GEN_365; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_367 = 7'h6f == predictor_idx_2[6:0] ? predictor_111 : _GEN_366; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_368 = 7'h70 == predictor_idx_2[6:0] ? predictor_112 : _GEN_367; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_369 = 7'h71 == predictor_idx_2[6:0] ? predictor_113 : _GEN_368; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_370 = 7'h72 == predictor_idx_2[6:0] ? predictor_114 : _GEN_369; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_371 = 7'h73 == predictor_idx_2[6:0] ? predictor_115 : _GEN_370; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_372 = 7'h74 == predictor_idx_2[6:0] ? predictor_116 : _GEN_371; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_373 = 7'h75 == predictor_idx_2[6:0] ? predictor_117 : _GEN_372; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_374 = 7'h76 == predictor_idx_2[6:0] ? predictor_118 : _GEN_373; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_375 = 7'h77 == predictor_idx_2[6:0] ? predictor_119 : _GEN_374; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_376 = 7'h78 == predictor_idx_2[6:0] ? predictor_120 : _GEN_375; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_377 = 7'h79 == predictor_idx_2[6:0] ? predictor_121 : _GEN_376; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_378 = 7'h7a == predictor_idx_2[6:0] ? predictor_122 : _GEN_377; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_379 = 7'h7b == predictor_idx_2[6:0] ? predictor_123 : _GEN_378; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_380 = 7'h7c == predictor_idx_2[6:0] ? predictor_124 : _GEN_379; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_381 = 7'h7d == predictor_idx_2[6:0] ? predictor_125 : _GEN_380; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_382 = 7'h7e == predictor_idx_2[6:0] ? predictor_126 : _GEN_381; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_383 = 7'h7f == predictor_idx_2[6:0] ? predictor_127 : _GEN_382; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire  predict_mask_2 = _GEN_383[1]; // @[Bpu.scala 96:62]
  wire [1:0] _GEN_385 = 7'h1 == predictor_idx_3[6:0] ? predictor_1 : predictor_0; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_386 = 7'h2 == predictor_idx_3[6:0] ? predictor_2 : _GEN_385; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_387 = 7'h3 == predictor_idx_3[6:0] ? predictor_3 : _GEN_386; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_388 = 7'h4 == predictor_idx_3[6:0] ? predictor_4 : _GEN_387; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_389 = 7'h5 == predictor_idx_3[6:0] ? predictor_5 : _GEN_388; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_390 = 7'h6 == predictor_idx_3[6:0] ? predictor_6 : _GEN_389; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_391 = 7'h7 == predictor_idx_3[6:0] ? predictor_7 : _GEN_390; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_392 = 7'h8 == predictor_idx_3[6:0] ? predictor_8 : _GEN_391; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_393 = 7'h9 == predictor_idx_3[6:0] ? predictor_9 : _GEN_392; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_394 = 7'ha == predictor_idx_3[6:0] ? predictor_10 : _GEN_393; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_395 = 7'hb == predictor_idx_3[6:0] ? predictor_11 : _GEN_394; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_396 = 7'hc == predictor_idx_3[6:0] ? predictor_12 : _GEN_395; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_397 = 7'hd == predictor_idx_3[6:0] ? predictor_13 : _GEN_396; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_398 = 7'he == predictor_idx_3[6:0] ? predictor_14 : _GEN_397; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_399 = 7'hf == predictor_idx_3[6:0] ? predictor_15 : _GEN_398; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_400 = 7'h10 == predictor_idx_3[6:0] ? predictor_16 : _GEN_399; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_401 = 7'h11 == predictor_idx_3[6:0] ? predictor_17 : _GEN_400; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_402 = 7'h12 == predictor_idx_3[6:0] ? predictor_18 : _GEN_401; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_403 = 7'h13 == predictor_idx_3[6:0] ? predictor_19 : _GEN_402; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_404 = 7'h14 == predictor_idx_3[6:0] ? predictor_20 : _GEN_403; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_405 = 7'h15 == predictor_idx_3[6:0] ? predictor_21 : _GEN_404; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_406 = 7'h16 == predictor_idx_3[6:0] ? predictor_22 : _GEN_405; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_407 = 7'h17 == predictor_idx_3[6:0] ? predictor_23 : _GEN_406; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_408 = 7'h18 == predictor_idx_3[6:0] ? predictor_24 : _GEN_407; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_409 = 7'h19 == predictor_idx_3[6:0] ? predictor_25 : _GEN_408; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_410 = 7'h1a == predictor_idx_3[6:0] ? predictor_26 : _GEN_409; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_411 = 7'h1b == predictor_idx_3[6:0] ? predictor_27 : _GEN_410; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_412 = 7'h1c == predictor_idx_3[6:0] ? predictor_28 : _GEN_411; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_413 = 7'h1d == predictor_idx_3[6:0] ? predictor_29 : _GEN_412; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_414 = 7'h1e == predictor_idx_3[6:0] ? predictor_30 : _GEN_413; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_415 = 7'h1f == predictor_idx_3[6:0] ? predictor_31 : _GEN_414; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_416 = 7'h20 == predictor_idx_3[6:0] ? predictor_32 : _GEN_415; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_417 = 7'h21 == predictor_idx_3[6:0] ? predictor_33 : _GEN_416; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_418 = 7'h22 == predictor_idx_3[6:0] ? predictor_34 : _GEN_417; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_419 = 7'h23 == predictor_idx_3[6:0] ? predictor_35 : _GEN_418; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_420 = 7'h24 == predictor_idx_3[6:0] ? predictor_36 : _GEN_419; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_421 = 7'h25 == predictor_idx_3[6:0] ? predictor_37 : _GEN_420; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_422 = 7'h26 == predictor_idx_3[6:0] ? predictor_38 : _GEN_421; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_423 = 7'h27 == predictor_idx_3[6:0] ? predictor_39 : _GEN_422; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_424 = 7'h28 == predictor_idx_3[6:0] ? predictor_40 : _GEN_423; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_425 = 7'h29 == predictor_idx_3[6:0] ? predictor_41 : _GEN_424; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_426 = 7'h2a == predictor_idx_3[6:0] ? predictor_42 : _GEN_425; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_427 = 7'h2b == predictor_idx_3[6:0] ? predictor_43 : _GEN_426; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_428 = 7'h2c == predictor_idx_3[6:0] ? predictor_44 : _GEN_427; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_429 = 7'h2d == predictor_idx_3[6:0] ? predictor_45 : _GEN_428; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_430 = 7'h2e == predictor_idx_3[6:0] ? predictor_46 : _GEN_429; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_431 = 7'h2f == predictor_idx_3[6:0] ? predictor_47 : _GEN_430; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_432 = 7'h30 == predictor_idx_3[6:0] ? predictor_48 : _GEN_431; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_433 = 7'h31 == predictor_idx_3[6:0] ? predictor_49 : _GEN_432; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_434 = 7'h32 == predictor_idx_3[6:0] ? predictor_50 : _GEN_433; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_435 = 7'h33 == predictor_idx_3[6:0] ? predictor_51 : _GEN_434; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_436 = 7'h34 == predictor_idx_3[6:0] ? predictor_52 : _GEN_435; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_437 = 7'h35 == predictor_idx_3[6:0] ? predictor_53 : _GEN_436; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_438 = 7'h36 == predictor_idx_3[6:0] ? predictor_54 : _GEN_437; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_439 = 7'h37 == predictor_idx_3[6:0] ? predictor_55 : _GEN_438; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_440 = 7'h38 == predictor_idx_3[6:0] ? predictor_56 : _GEN_439; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_441 = 7'h39 == predictor_idx_3[6:0] ? predictor_57 : _GEN_440; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_442 = 7'h3a == predictor_idx_3[6:0] ? predictor_58 : _GEN_441; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_443 = 7'h3b == predictor_idx_3[6:0] ? predictor_59 : _GEN_442; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_444 = 7'h3c == predictor_idx_3[6:0] ? predictor_60 : _GEN_443; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_445 = 7'h3d == predictor_idx_3[6:0] ? predictor_61 : _GEN_444; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_446 = 7'h3e == predictor_idx_3[6:0] ? predictor_62 : _GEN_445; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_447 = 7'h3f == predictor_idx_3[6:0] ? predictor_63 : _GEN_446; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_448 = 7'h40 == predictor_idx_3[6:0] ? predictor_64 : _GEN_447; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_449 = 7'h41 == predictor_idx_3[6:0] ? predictor_65 : _GEN_448; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_450 = 7'h42 == predictor_idx_3[6:0] ? predictor_66 : _GEN_449; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_451 = 7'h43 == predictor_idx_3[6:0] ? predictor_67 : _GEN_450; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_452 = 7'h44 == predictor_idx_3[6:0] ? predictor_68 : _GEN_451; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_453 = 7'h45 == predictor_idx_3[6:0] ? predictor_69 : _GEN_452; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_454 = 7'h46 == predictor_idx_3[6:0] ? predictor_70 : _GEN_453; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_455 = 7'h47 == predictor_idx_3[6:0] ? predictor_71 : _GEN_454; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_456 = 7'h48 == predictor_idx_3[6:0] ? predictor_72 : _GEN_455; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_457 = 7'h49 == predictor_idx_3[6:0] ? predictor_73 : _GEN_456; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_458 = 7'h4a == predictor_idx_3[6:0] ? predictor_74 : _GEN_457; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_459 = 7'h4b == predictor_idx_3[6:0] ? predictor_75 : _GEN_458; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_460 = 7'h4c == predictor_idx_3[6:0] ? predictor_76 : _GEN_459; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_461 = 7'h4d == predictor_idx_3[6:0] ? predictor_77 : _GEN_460; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_462 = 7'h4e == predictor_idx_3[6:0] ? predictor_78 : _GEN_461; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_463 = 7'h4f == predictor_idx_3[6:0] ? predictor_79 : _GEN_462; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_464 = 7'h50 == predictor_idx_3[6:0] ? predictor_80 : _GEN_463; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_465 = 7'h51 == predictor_idx_3[6:0] ? predictor_81 : _GEN_464; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_466 = 7'h52 == predictor_idx_3[6:0] ? predictor_82 : _GEN_465; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_467 = 7'h53 == predictor_idx_3[6:0] ? predictor_83 : _GEN_466; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_468 = 7'h54 == predictor_idx_3[6:0] ? predictor_84 : _GEN_467; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_469 = 7'h55 == predictor_idx_3[6:0] ? predictor_85 : _GEN_468; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_470 = 7'h56 == predictor_idx_3[6:0] ? predictor_86 : _GEN_469; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_471 = 7'h57 == predictor_idx_3[6:0] ? predictor_87 : _GEN_470; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_472 = 7'h58 == predictor_idx_3[6:0] ? predictor_88 : _GEN_471; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_473 = 7'h59 == predictor_idx_3[6:0] ? predictor_89 : _GEN_472; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_474 = 7'h5a == predictor_idx_3[6:0] ? predictor_90 : _GEN_473; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_475 = 7'h5b == predictor_idx_3[6:0] ? predictor_91 : _GEN_474; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_476 = 7'h5c == predictor_idx_3[6:0] ? predictor_92 : _GEN_475; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_477 = 7'h5d == predictor_idx_3[6:0] ? predictor_93 : _GEN_476; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_478 = 7'h5e == predictor_idx_3[6:0] ? predictor_94 : _GEN_477; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_479 = 7'h5f == predictor_idx_3[6:0] ? predictor_95 : _GEN_478; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_480 = 7'h60 == predictor_idx_3[6:0] ? predictor_96 : _GEN_479; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_481 = 7'h61 == predictor_idx_3[6:0] ? predictor_97 : _GEN_480; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_482 = 7'h62 == predictor_idx_3[6:0] ? predictor_98 : _GEN_481; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_483 = 7'h63 == predictor_idx_3[6:0] ? predictor_99 : _GEN_482; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_484 = 7'h64 == predictor_idx_3[6:0] ? predictor_100 : _GEN_483; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_485 = 7'h65 == predictor_idx_3[6:0] ? predictor_101 : _GEN_484; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_486 = 7'h66 == predictor_idx_3[6:0] ? predictor_102 : _GEN_485; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_487 = 7'h67 == predictor_idx_3[6:0] ? predictor_103 : _GEN_486; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_488 = 7'h68 == predictor_idx_3[6:0] ? predictor_104 : _GEN_487; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_489 = 7'h69 == predictor_idx_3[6:0] ? predictor_105 : _GEN_488; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_490 = 7'h6a == predictor_idx_3[6:0] ? predictor_106 : _GEN_489; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_491 = 7'h6b == predictor_idx_3[6:0] ? predictor_107 : _GEN_490; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_492 = 7'h6c == predictor_idx_3[6:0] ? predictor_108 : _GEN_491; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_493 = 7'h6d == predictor_idx_3[6:0] ? predictor_109 : _GEN_492; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_494 = 7'h6e == predictor_idx_3[6:0] ? predictor_110 : _GEN_493; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_495 = 7'h6f == predictor_idx_3[6:0] ? predictor_111 : _GEN_494; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_496 = 7'h70 == predictor_idx_3[6:0] ? predictor_112 : _GEN_495; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_497 = 7'h71 == predictor_idx_3[6:0] ? predictor_113 : _GEN_496; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_498 = 7'h72 == predictor_idx_3[6:0] ? predictor_114 : _GEN_497; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_499 = 7'h73 == predictor_idx_3[6:0] ? predictor_115 : _GEN_498; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_500 = 7'h74 == predictor_idx_3[6:0] ? predictor_116 : _GEN_499; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_501 = 7'h75 == predictor_idx_3[6:0] ? predictor_117 : _GEN_500; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_502 = 7'h76 == predictor_idx_3[6:0] ? predictor_118 : _GEN_501; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_503 = 7'h77 == predictor_idx_3[6:0] ? predictor_119 : _GEN_502; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_504 = 7'h78 == predictor_idx_3[6:0] ? predictor_120 : _GEN_503; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_505 = 7'h79 == predictor_idx_3[6:0] ? predictor_121 : _GEN_504; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_506 = 7'h7a == predictor_idx_3[6:0] ? predictor_122 : _GEN_505; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_507 = 7'h7b == predictor_idx_3[6:0] ? predictor_123 : _GEN_506; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_508 = 7'h7c == predictor_idx_3[6:0] ? predictor_124 : _GEN_507; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_509 = 7'h7d == predictor_idx_3[6:0] ? predictor_125 : _GEN_508; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_510 = 7'h7e == predictor_idx_3[6:0] ? predictor_126 : _GEN_509; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_511 = 7'h7f == predictor_idx_3[6:0] ? predictor_127 : _GEN_510; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire  predict_mask_3 = _GEN_511[1]; // @[Bpu.scala 96:62]
  wire [1:0] _GEN_513 = 7'h1 == predictor_idx_4[6:0] ? predictor_1 : predictor_0; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_514 = 7'h2 == predictor_idx_4[6:0] ? predictor_2 : _GEN_513; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_515 = 7'h3 == predictor_idx_4[6:0] ? predictor_3 : _GEN_514; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_516 = 7'h4 == predictor_idx_4[6:0] ? predictor_4 : _GEN_515; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_517 = 7'h5 == predictor_idx_4[6:0] ? predictor_5 : _GEN_516; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_518 = 7'h6 == predictor_idx_4[6:0] ? predictor_6 : _GEN_517; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_519 = 7'h7 == predictor_idx_4[6:0] ? predictor_7 : _GEN_518; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_520 = 7'h8 == predictor_idx_4[6:0] ? predictor_8 : _GEN_519; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_521 = 7'h9 == predictor_idx_4[6:0] ? predictor_9 : _GEN_520; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_522 = 7'ha == predictor_idx_4[6:0] ? predictor_10 : _GEN_521; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_523 = 7'hb == predictor_idx_4[6:0] ? predictor_11 : _GEN_522; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_524 = 7'hc == predictor_idx_4[6:0] ? predictor_12 : _GEN_523; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_525 = 7'hd == predictor_idx_4[6:0] ? predictor_13 : _GEN_524; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_526 = 7'he == predictor_idx_4[6:0] ? predictor_14 : _GEN_525; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_527 = 7'hf == predictor_idx_4[6:0] ? predictor_15 : _GEN_526; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_528 = 7'h10 == predictor_idx_4[6:0] ? predictor_16 : _GEN_527; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_529 = 7'h11 == predictor_idx_4[6:0] ? predictor_17 : _GEN_528; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_530 = 7'h12 == predictor_idx_4[6:0] ? predictor_18 : _GEN_529; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_531 = 7'h13 == predictor_idx_4[6:0] ? predictor_19 : _GEN_530; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_532 = 7'h14 == predictor_idx_4[6:0] ? predictor_20 : _GEN_531; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_533 = 7'h15 == predictor_idx_4[6:0] ? predictor_21 : _GEN_532; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_534 = 7'h16 == predictor_idx_4[6:0] ? predictor_22 : _GEN_533; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_535 = 7'h17 == predictor_idx_4[6:0] ? predictor_23 : _GEN_534; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_536 = 7'h18 == predictor_idx_4[6:0] ? predictor_24 : _GEN_535; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_537 = 7'h19 == predictor_idx_4[6:0] ? predictor_25 : _GEN_536; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_538 = 7'h1a == predictor_idx_4[6:0] ? predictor_26 : _GEN_537; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_539 = 7'h1b == predictor_idx_4[6:0] ? predictor_27 : _GEN_538; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_540 = 7'h1c == predictor_idx_4[6:0] ? predictor_28 : _GEN_539; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_541 = 7'h1d == predictor_idx_4[6:0] ? predictor_29 : _GEN_540; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_542 = 7'h1e == predictor_idx_4[6:0] ? predictor_30 : _GEN_541; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_543 = 7'h1f == predictor_idx_4[6:0] ? predictor_31 : _GEN_542; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_544 = 7'h20 == predictor_idx_4[6:0] ? predictor_32 : _GEN_543; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_545 = 7'h21 == predictor_idx_4[6:0] ? predictor_33 : _GEN_544; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_546 = 7'h22 == predictor_idx_4[6:0] ? predictor_34 : _GEN_545; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_547 = 7'h23 == predictor_idx_4[6:0] ? predictor_35 : _GEN_546; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_548 = 7'h24 == predictor_idx_4[6:0] ? predictor_36 : _GEN_547; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_549 = 7'h25 == predictor_idx_4[6:0] ? predictor_37 : _GEN_548; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_550 = 7'h26 == predictor_idx_4[6:0] ? predictor_38 : _GEN_549; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_551 = 7'h27 == predictor_idx_4[6:0] ? predictor_39 : _GEN_550; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_552 = 7'h28 == predictor_idx_4[6:0] ? predictor_40 : _GEN_551; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_553 = 7'h29 == predictor_idx_4[6:0] ? predictor_41 : _GEN_552; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_554 = 7'h2a == predictor_idx_4[6:0] ? predictor_42 : _GEN_553; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_555 = 7'h2b == predictor_idx_4[6:0] ? predictor_43 : _GEN_554; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_556 = 7'h2c == predictor_idx_4[6:0] ? predictor_44 : _GEN_555; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_557 = 7'h2d == predictor_idx_4[6:0] ? predictor_45 : _GEN_556; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_558 = 7'h2e == predictor_idx_4[6:0] ? predictor_46 : _GEN_557; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_559 = 7'h2f == predictor_idx_4[6:0] ? predictor_47 : _GEN_558; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_560 = 7'h30 == predictor_idx_4[6:0] ? predictor_48 : _GEN_559; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_561 = 7'h31 == predictor_idx_4[6:0] ? predictor_49 : _GEN_560; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_562 = 7'h32 == predictor_idx_4[6:0] ? predictor_50 : _GEN_561; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_563 = 7'h33 == predictor_idx_4[6:0] ? predictor_51 : _GEN_562; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_564 = 7'h34 == predictor_idx_4[6:0] ? predictor_52 : _GEN_563; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_565 = 7'h35 == predictor_idx_4[6:0] ? predictor_53 : _GEN_564; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_566 = 7'h36 == predictor_idx_4[6:0] ? predictor_54 : _GEN_565; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_567 = 7'h37 == predictor_idx_4[6:0] ? predictor_55 : _GEN_566; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_568 = 7'h38 == predictor_idx_4[6:0] ? predictor_56 : _GEN_567; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_569 = 7'h39 == predictor_idx_4[6:0] ? predictor_57 : _GEN_568; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_570 = 7'h3a == predictor_idx_4[6:0] ? predictor_58 : _GEN_569; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_571 = 7'h3b == predictor_idx_4[6:0] ? predictor_59 : _GEN_570; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_572 = 7'h3c == predictor_idx_4[6:0] ? predictor_60 : _GEN_571; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_573 = 7'h3d == predictor_idx_4[6:0] ? predictor_61 : _GEN_572; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_574 = 7'h3e == predictor_idx_4[6:0] ? predictor_62 : _GEN_573; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_575 = 7'h3f == predictor_idx_4[6:0] ? predictor_63 : _GEN_574; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_576 = 7'h40 == predictor_idx_4[6:0] ? predictor_64 : _GEN_575; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_577 = 7'h41 == predictor_idx_4[6:0] ? predictor_65 : _GEN_576; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_578 = 7'h42 == predictor_idx_4[6:0] ? predictor_66 : _GEN_577; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_579 = 7'h43 == predictor_idx_4[6:0] ? predictor_67 : _GEN_578; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_580 = 7'h44 == predictor_idx_4[6:0] ? predictor_68 : _GEN_579; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_581 = 7'h45 == predictor_idx_4[6:0] ? predictor_69 : _GEN_580; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_582 = 7'h46 == predictor_idx_4[6:0] ? predictor_70 : _GEN_581; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_583 = 7'h47 == predictor_idx_4[6:0] ? predictor_71 : _GEN_582; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_584 = 7'h48 == predictor_idx_4[6:0] ? predictor_72 : _GEN_583; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_585 = 7'h49 == predictor_idx_4[6:0] ? predictor_73 : _GEN_584; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_586 = 7'h4a == predictor_idx_4[6:0] ? predictor_74 : _GEN_585; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_587 = 7'h4b == predictor_idx_4[6:0] ? predictor_75 : _GEN_586; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_588 = 7'h4c == predictor_idx_4[6:0] ? predictor_76 : _GEN_587; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_589 = 7'h4d == predictor_idx_4[6:0] ? predictor_77 : _GEN_588; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_590 = 7'h4e == predictor_idx_4[6:0] ? predictor_78 : _GEN_589; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_591 = 7'h4f == predictor_idx_4[6:0] ? predictor_79 : _GEN_590; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_592 = 7'h50 == predictor_idx_4[6:0] ? predictor_80 : _GEN_591; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_593 = 7'h51 == predictor_idx_4[6:0] ? predictor_81 : _GEN_592; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_594 = 7'h52 == predictor_idx_4[6:0] ? predictor_82 : _GEN_593; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_595 = 7'h53 == predictor_idx_4[6:0] ? predictor_83 : _GEN_594; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_596 = 7'h54 == predictor_idx_4[6:0] ? predictor_84 : _GEN_595; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_597 = 7'h55 == predictor_idx_4[6:0] ? predictor_85 : _GEN_596; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_598 = 7'h56 == predictor_idx_4[6:0] ? predictor_86 : _GEN_597; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_599 = 7'h57 == predictor_idx_4[6:0] ? predictor_87 : _GEN_598; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_600 = 7'h58 == predictor_idx_4[6:0] ? predictor_88 : _GEN_599; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_601 = 7'h59 == predictor_idx_4[6:0] ? predictor_89 : _GEN_600; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_602 = 7'h5a == predictor_idx_4[6:0] ? predictor_90 : _GEN_601; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_603 = 7'h5b == predictor_idx_4[6:0] ? predictor_91 : _GEN_602; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_604 = 7'h5c == predictor_idx_4[6:0] ? predictor_92 : _GEN_603; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_605 = 7'h5d == predictor_idx_4[6:0] ? predictor_93 : _GEN_604; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_606 = 7'h5e == predictor_idx_4[6:0] ? predictor_94 : _GEN_605; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_607 = 7'h5f == predictor_idx_4[6:0] ? predictor_95 : _GEN_606; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_608 = 7'h60 == predictor_idx_4[6:0] ? predictor_96 : _GEN_607; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_609 = 7'h61 == predictor_idx_4[6:0] ? predictor_97 : _GEN_608; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_610 = 7'h62 == predictor_idx_4[6:0] ? predictor_98 : _GEN_609; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_611 = 7'h63 == predictor_idx_4[6:0] ? predictor_99 : _GEN_610; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_612 = 7'h64 == predictor_idx_4[6:0] ? predictor_100 : _GEN_611; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_613 = 7'h65 == predictor_idx_4[6:0] ? predictor_101 : _GEN_612; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_614 = 7'h66 == predictor_idx_4[6:0] ? predictor_102 : _GEN_613; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_615 = 7'h67 == predictor_idx_4[6:0] ? predictor_103 : _GEN_614; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_616 = 7'h68 == predictor_idx_4[6:0] ? predictor_104 : _GEN_615; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_617 = 7'h69 == predictor_idx_4[6:0] ? predictor_105 : _GEN_616; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_618 = 7'h6a == predictor_idx_4[6:0] ? predictor_106 : _GEN_617; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_619 = 7'h6b == predictor_idx_4[6:0] ? predictor_107 : _GEN_618; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_620 = 7'h6c == predictor_idx_4[6:0] ? predictor_108 : _GEN_619; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_621 = 7'h6d == predictor_idx_4[6:0] ? predictor_109 : _GEN_620; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_622 = 7'h6e == predictor_idx_4[6:0] ? predictor_110 : _GEN_621; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_623 = 7'h6f == predictor_idx_4[6:0] ? predictor_111 : _GEN_622; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_624 = 7'h70 == predictor_idx_4[6:0] ? predictor_112 : _GEN_623; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_625 = 7'h71 == predictor_idx_4[6:0] ? predictor_113 : _GEN_624; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_626 = 7'h72 == predictor_idx_4[6:0] ? predictor_114 : _GEN_625; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_627 = 7'h73 == predictor_idx_4[6:0] ? predictor_115 : _GEN_626; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_628 = 7'h74 == predictor_idx_4[6:0] ? predictor_116 : _GEN_627; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_629 = 7'h75 == predictor_idx_4[6:0] ? predictor_117 : _GEN_628; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_630 = 7'h76 == predictor_idx_4[6:0] ? predictor_118 : _GEN_629; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_631 = 7'h77 == predictor_idx_4[6:0] ? predictor_119 : _GEN_630; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_632 = 7'h78 == predictor_idx_4[6:0] ? predictor_120 : _GEN_631; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_633 = 7'h79 == predictor_idx_4[6:0] ? predictor_121 : _GEN_632; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_634 = 7'h7a == predictor_idx_4[6:0] ? predictor_122 : _GEN_633; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_635 = 7'h7b == predictor_idx_4[6:0] ? predictor_123 : _GEN_634; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_636 = 7'h7c == predictor_idx_4[6:0] ? predictor_124 : _GEN_635; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_637 = 7'h7d == predictor_idx_4[6:0] ? predictor_125 : _GEN_636; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_638 = 7'h7e == predictor_idx_4[6:0] ? predictor_126 : _GEN_637; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_639 = 7'h7f == predictor_idx_4[6:0] ? predictor_127 : _GEN_638; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire  predict_mask_4 = _GEN_639[1]; // @[Bpu.scala 96:62]
  wire [1:0] _GEN_641 = 7'h1 == predictor_idx_5[6:0] ? predictor_1 : predictor_0; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_642 = 7'h2 == predictor_idx_5[6:0] ? predictor_2 : _GEN_641; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_643 = 7'h3 == predictor_idx_5[6:0] ? predictor_3 : _GEN_642; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_644 = 7'h4 == predictor_idx_5[6:0] ? predictor_4 : _GEN_643; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_645 = 7'h5 == predictor_idx_5[6:0] ? predictor_5 : _GEN_644; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_646 = 7'h6 == predictor_idx_5[6:0] ? predictor_6 : _GEN_645; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_647 = 7'h7 == predictor_idx_5[6:0] ? predictor_7 : _GEN_646; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_648 = 7'h8 == predictor_idx_5[6:0] ? predictor_8 : _GEN_647; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_649 = 7'h9 == predictor_idx_5[6:0] ? predictor_9 : _GEN_648; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_650 = 7'ha == predictor_idx_5[6:0] ? predictor_10 : _GEN_649; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_651 = 7'hb == predictor_idx_5[6:0] ? predictor_11 : _GEN_650; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_652 = 7'hc == predictor_idx_5[6:0] ? predictor_12 : _GEN_651; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_653 = 7'hd == predictor_idx_5[6:0] ? predictor_13 : _GEN_652; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_654 = 7'he == predictor_idx_5[6:0] ? predictor_14 : _GEN_653; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_655 = 7'hf == predictor_idx_5[6:0] ? predictor_15 : _GEN_654; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_656 = 7'h10 == predictor_idx_5[6:0] ? predictor_16 : _GEN_655; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_657 = 7'h11 == predictor_idx_5[6:0] ? predictor_17 : _GEN_656; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_658 = 7'h12 == predictor_idx_5[6:0] ? predictor_18 : _GEN_657; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_659 = 7'h13 == predictor_idx_5[6:0] ? predictor_19 : _GEN_658; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_660 = 7'h14 == predictor_idx_5[6:0] ? predictor_20 : _GEN_659; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_661 = 7'h15 == predictor_idx_5[6:0] ? predictor_21 : _GEN_660; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_662 = 7'h16 == predictor_idx_5[6:0] ? predictor_22 : _GEN_661; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_663 = 7'h17 == predictor_idx_5[6:0] ? predictor_23 : _GEN_662; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_664 = 7'h18 == predictor_idx_5[6:0] ? predictor_24 : _GEN_663; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_665 = 7'h19 == predictor_idx_5[6:0] ? predictor_25 : _GEN_664; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_666 = 7'h1a == predictor_idx_5[6:0] ? predictor_26 : _GEN_665; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_667 = 7'h1b == predictor_idx_5[6:0] ? predictor_27 : _GEN_666; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_668 = 7'h1c == predictor_idx_5[6:0] ? predictor_28 : _GEN_667; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_669 = 7'h1d == predictor_idx_5[6:0] ? predictor_29 : _GEN_668; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_670 = 7'h1e == predictor_idx_5[6:0] ? predictor_30 : _GEN_669; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_671 = 7'h1f == predictor_idx_5[6:0] ? predictor_31 : _GEN_670; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_672 = 7'h20 == predictor_idx_5[6:0] ? predictor_32 : _GEN_671; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_673 = 7'h21 == predictor_idx_5[6:0] ? predictor_33 : _GEN_672; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_674 = 7'h22 == predictor_idx_5[6:0] ? predictor_34 : _GEN_673; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_675 = 7'h23 == predictor_idx_5[6:0] ? predictor_35 : _GEN_674; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_676 = 7'h24 == predictor_idx_5[6:0] ? predictor_36 : _GEN_675; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_677 = 7'h25 == predictor_idx_5[6:0] ? predictor_37 : _GEN_676; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_678 = 7'h26 == predictor_idx_5[6:0] ? predictor_38 : _GEN_677; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_679 = 7'h27 == predictor_idx_5[6:0] ? predictor_39 : _GEN_678; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_680 = 7'h28 == predictor_idx_5[6:0] ? predictor_40 : _GEN_679; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_681 = 7'h29 == predictor_idx_5[6:0] ? predictor_41 : _GEN_680; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_682 = 7'h2a == predictor_idx_5[6:0] ? predictor_42 : _GEN_681; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_683 = 7'h2b == predictor_idx_5[6:0] ? predictor_43 : _GEN_682; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_684 = 7'h2c == predictor_idx_5[6:0] ? predictor_44 : _GEN_683; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_685 = 7'h2d == predictor_idx_5[6:0] ? predictor_45 : _GEN_684; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_686 = 7'h2e == predictor_idx_5[6:0] ? predictor_46 : _GEN_685; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_687 = 7'h2f == predictor_idx_5[6:0] ? predictor_47 : _GEN_686; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_688 = 7'h30 == predictor_idx_5[6:0] ? predictor_48 : _GEN_687; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_689 = 7'h31 == predictor_idx_5[6:0] ? predictor_49 : _GEN_688; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_690 = 7'h32 == predictor_idx_5[6:0] ? predictor_50 : _GEN_689; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_691 = 7'h33 == predictor_idx_5[6:0] ? predictor_51 : _GEN_690; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_692 = 7'h34 == predictor_idx_5[6:0] ? predictor_52 : _GEN_691; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_693 = 7'h35 == predictor_idx_5[6:0] ? predictor_53 : _GEN_692; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_694 = 7'h36 == predictor_idx_5[6:0] ? predictor_54 : _GEN_693; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_695 = 7'h37 == predictor_idx_5[6:0] ? predictor_55 : _GEN_694; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_696 = 7'h38 == predictor_idx_5[6:0] ? predictor_56 : _GEN_695; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_697 = 7'h39 == predictor_idx_5[6:0] ? predictor_57 : _GEN_696; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_698 = 7'h3a == predictor_idx_5[6:0] ? predictor_58 : _GEN_697; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_699 = 7'h3b == predictor_idx_5[6:0] ? predictor_59 : _GEN_698; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_700 = 7'h3c == predictor_idx_5[6:0] ? predictor_60 : _GEN_699; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_701 = 7'h3d == predictor_idx_5[6:0] ? predictor_61 : _GEN_700; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_702 = 7'h3e == predictor_idx_5[6:0] ? predictor_62 : _GEN_701; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_703 = 7'h3f == predictor_idx_5[6:0] ? predictor_63 : _GEN_702; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_704 = 7'h40 == predictor_idx_5[6:0] ? predictor_64 : _GEN_703; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_705 = 7'h41 == predictor_idx_5[6:0] ? predictor_65 : _GEN_704; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_706 = 7'h42 == predictor_idx_5[6:0] ? predictor_66 : _GEN_705; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_707 = 7'h43 == predictor_idx_5[6:0] ? predictor_67 : _GEN_706; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_708 = 7'h44 == predictor_idx_5[6:0] ? predictor_68 : _GEN_707; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_709 = 7'h45 == predictor_idx_5[6:0] ? predictor_69 : _GEN_708; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_710 = 7'h46 == predictor_idx_5[6:0] ? predictor_70 : _GEN_709; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_711 = 7'h47 == predictor_idx_5[6:0] ? predictor_71 : _GEN_710; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_712 = 7'h48 == predictor_idx_5[6:0] ? predictor_72 : _GEN_711; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_713 = 7'h49 == predictor_idx_5[6:0] ? predictor_73 : _GEN_712; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_714 = 7'h4a == predictor_idx_5[6:0] ? predictor_74 : _GEN_713; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_715 = 7'h4b == predictor_idx_5[6:0] ? predictor_75 : _GEN_714; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_716 = 7'h4c == predictor_idx_5[6:0] ? predictor_76 : _GEN_715; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_717 = 7'h4d == predictor_idx_5[6:0] ? predictor_77 : _GEN_716; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_718 = 7'h4e == predictor_idx_5[6:0] ? predictor_78 : _GEN_717; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_719 = 7'h4f == predictor_idx_5[6:0] ? predictor_79 : _GEN_718; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_720 = 7'h50 == predictor_idx_5[6:0] ? predictor_80 : _GEN_719; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_721 = 7'h51 == predictor_idx_5[6:0] ? predictor_81 : _GEN_720; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_722 = 7'h52 == predictor_idx_5[6:0] ? predictor_82 : _GEN_721; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_723 = 7'h53 == predictor_idx_5[6:0] ? predictor_83 : _GEN_722; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_724 = 7'h54 == predictor_idx_5[6:0] ? predictor_84 : _GEN_723; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_725 = 7'h55 == predictor_idx_5[6:0] ? predictor_85 : _GEN_724; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_726 = 7'h56 == predictor_idx_5[6:0] ? predictor_86 : _GEN_725; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_727 = 7'h57 == predictor_idx_5[6:0] ? predictor_87 : _GEN_726; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_728 = 7'h58 == predictor_idx_5[6:0] ? predictor_88 : _GEN_727; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_729 = 7'h59 == predictor_idx_5[6:0] ? predictor_89 : _GEN_728; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_730 = 7'h5a == predictor_idx_5[6:0] ? predictor_90 : _GEN_729; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_731 = 7'h5b == predictor_idx_5[6:0] ? predictor_91 : _GEN_730; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_732 = 7'h5c == predictor_idx_5[6:0] ? predictor_92 : _GEN_731; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_733 = 7'h5d == predictor_idx_5[6:0] ? predictor_93 : _GEN_732; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_734 = 7'h5e == predictor_idx_5[6:0] ? predictor_94 : _GEN_733; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_735 = 7'h5f == predictor_idx_5[6:0] ? predictor_95 : _GEN_734; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_736 = 7'h60 == predictor_idx_5[6:0] ? predictor_96 : _GEN_735; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_737 = 7'h61 == predictor_idx_5[6:0] ? predictor_97 : _GEN_736; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_738 = 7'h62 == predictor_idx_5[6:0] ? predictor_98 : _GEN_737; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_739 = 7'h63 == predictor_idx_5[6:0] ? predictor_99 : _GEN_738; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_740 = 7'h64 == predictor_idx_5[6:0] ? predictor_100 : _GEN_739; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_741 = 7'h65 == predictor_idx_5[6:0] ? predictor_101 : _GEN_740; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_742 = 7'h66 == predictor_idx_5[6:0] ? predictor_102 : _GEN_741; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_743 = 7'h67 == predictor_idx_5[6:0] ? predictor_103 : _GEN_742; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_744 = 7'h68 == predictor_idx_5[6:0] ? predictor_104 : _GEN_743; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_745 = 7'h69 == predictor_idx_5[6:0] ? predictor_105 : _GEN_744; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_746 = 7'h6a == predictor_idx_5[6:0] ? predictor_106 : _GEN_745; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_747 = 7'h6b == predictor_idx_5[6:0] ? predictor_107 : _GEN_746; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_748 = 7'h6c == predictor_idx_5[6:0] ? predictor_108 : _GEN_747; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_749 = 7'h6d == predictor_idx_5[6:0] ? predictor_109 : _GEN_748; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_750 = 7'h6e == predictor_idx_5[6:0] ? predictor_110 : _GEN_749; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_751 = 7'h6f == predictor_idx_5[6:0] ? predictor_111 : _GEN_750; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_752 = 7'h70 == predictor_idx_5[6:0] ? predictor_112 : _GEN_751; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_753 = 7'h71 == predictor_idx_5[6:0] ? predictor_113 : _GEN_752; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_754 = 7'h72 == predictor_idx_5[6:0] ? predictor_114 : _GEN_753; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_755 = 7'h73 == predictor_idx_5[6:0] ? predictor_115 : _GEN_754; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_756 = 7'h74 == predictor_idx_5[6:0] ? predictor_116 : _GEN_755; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_757 = 7'h75 == predictor_idx_5[6:0] ? predictor_117 : _GEN_756; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_758 = 7'h76 == predictor_idx_5[6:0] ? predictor_118 : _GEN_757; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_759 = 7'h77 == predictor_idx_5[6:0] ? predictor_119 : _GEN_758; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_760 = 7'h78 == predictor_idx_5[6:0] ? predictor_120 : _GEN_759; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_761 = 7'h79 == predictor_idx_5[6:0] ? predictor_121 : _GEN_760; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_762 = 7'h7a == predictor_idx_5[6:0] ? predictor_122 : _GEN_761; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_763 = 7'h7b == predictor_idx_5[6:0] ? predictor_123 : _GEN_762; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_764 = 7'h7c == predictor_idx_5[6:0] ? predictor_124 : _GEN_763; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_765 = 7'h7d == predictor_idx_5[6:0] ? predictor_125 : _GEN_764; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_766 = 7'h7e == predictor_idx_5[6:0] ? predictor_126 : _GEN_765; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_767 = 7'h7f == predictor_idx_5[6:0] ? predictor_127 : _GEN_766; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire  predict_mask_5 = _GEN_767[1]; // @[Bpu.scala 96:62]
  wire [1:0] _GEN_769 = 7'h1 == predictor_idx_6[6:0] ? predictor_1 : predictor_0; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_770 = 7'h2 == predictor_idx_6[6:0] ? predictor_2 : _GEN_769; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_771 = 7'h3 == predictor_idx_6[6:0] ? predictor_3 : _GEN_770; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_772 = 7'h4 == predictor_idx_6[6:0] ? predictor_4 : _GEN_771; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_773 = 7'h5 == predictor_idx_6[6:0] ? predictor_5 : _GEN_772; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_774 = 7'h6 == predictor_idx_6[6:0] ? predictor_6 : _GEN_773; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_775 = 7'h7 == predictor_idx_6[6:0] ? predictor_7 : _GEN_774; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_776 = 7'h8 == predictor_idx_6[6:0] ? predictor_8 : _GEN_775; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_777 = 7'h9 == predictor_idx_6[6:0] ? predictor_9 : _GEN_776; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_778 = 7'ha == predictor_idx_6[6:0] ? predictor_10 : _GEN_777; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_779 = 7'hb == predictor_idx_6[6:0] ? predictor_11 : _GEN_778; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_780 = 7'hc == predictor_idx_6[6:0] ? predictor_12 : _GEN_779; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_781 = 7'hd == predictor_idx_6[6:0] ? predictor_13 : _GEN_780; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_782 = 7'he == predictor_idx_6[6:0] ? predictor_14 : _GEN_781; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_783 = 7'hf == predictor_idx_6[6:0] ? predictor_15 : _GEN_782; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_784 = 7'h10 == predictor_idx_6[6:0] ? predictor_16 : _GEN_783; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_785 = 7'h11 == predictor_idx_6[6:0] ? predictor_17 : _GEN_784; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_786 = 7'h12 == predictor_idx_6[6:0] ? predictor_18 : _GEN_785; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_787 = 7'h13 == predictor_idx_6[6:0] ? predictor_19 : _GEN_786; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_788 = 7'h14 == predictor_idx_6[6:0] ? predictor_20 : _GEN_787; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_789 = 7'h15 == predictor_idx_6[6:0] ? predictor_21 : _GEN_788; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_790 = 7'h16 == predictor_idx_6[6:0] ? predictor_22 : _GEN_789; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_791 = 7'h17 == predictor_idx_6[6:0] ? predictor_23 : _GEN_790; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_792 = 7'h18 == predictor_idx_6[6:0] ? predictor_24 : _GEN_791; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_793 = 7'h19 == predictor_idx_6[6:0] ? predictor_25 : _GEN_792; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_794 = 7'h1a == predictor_idx_6[6:0] ? predictor_26 : _GEN_793; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_795 = 7'h1b == predictor_idx_6[6:0] ? predictor_27 : _GEN_794; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_796 = 7'h1c == predictor_idx_6[6:0] ? predictor_28 : _GEN_795; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_797 = 7'h1d == predictor_idx_6[6:0] ? predictor_29 : _GEN_796; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_798 = 7'h1e == predictor_idx_6[6:0] ? predictor_30 : _GEN_797; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_799 = 7'h1f == predictor_idx_6[6:0] ? predictor_31 : _GEN_798; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_800 = 7'h20 == predictor_idx_6[6:0] ? predictor_32 : _GEN_799; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_801 = 7'h21 == predictor_idx_6[6:0] ? predictor_33 : _GEN_800; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_802 = 7'h22 == predictor_idx_6[6:0] ? predictor_34 : _GEN_801; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_803 = 7'h23 == predictor_idx_6[6:0] ? predictor_35 : _GEN_802; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_804 = 7'h24 == predictor_idx_6[6:0] ? predictor_36 : _GEN_803; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_805 = 7'h25 == predictor_idx_6[6:0] ? predictor_37 : _GEN_804; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_806 = 7'h26 == predictor_idx_6[6:0] ? predictor_38 : _GEN_805; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_807 = 7'h27 == predictor_idx_6[6:0] ? predictor_39 : _GEN_806; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_808 = 7'h28 == predictor_idx_6[6:0] ? predictor_40 : _GEN_807; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_809 = 7'h29 == predictor_idx_6[6:0] ? predictor_41 : _GEN_808; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_810 = 7'h2a == predictor_idx_6[6:0] ? predictor_42 : _GEN_809; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_811 = 7'h2b == predictor_idx_6[6:0] ? predictor_43 : _GEN_810; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_812 = 7'h2c == predictor_idx_6[6:0] ? predictor_44 : _GEN_811; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_813 = 7'h2d == predictor_idx_6[6:0] ? predictor_45 : _GEN_812; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_814 = 7'h2e == predictor_idx_6[6:0] ? predictor_46 : _GEN_813; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_815 = 7'h2f == predictor_idx_6[6:0] ? predictor_47 : _GEN_814; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_816 = 7'h30 == predictor_idx_6[6:0] ? predictor_48 : _GEN_815; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_817 = 7'h31 == predictor_idx_6[6:0] ? predictor_49 : _GEN_816; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_818 = 7'h32 == predictor_idx_6[6:0] ? predictor_50 : _GEN_817; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_819 = 7'h33 == predictor_idx_6[6:0] ? predictor_51 : _GEN_818; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_820 = 7'h34 == predictor_idx_6[6:0] ? predictor_52 : _GEN_819; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_821 = 7'h35 == predictor_idx_6[6:0] ? predictor_53 : _GEN_820; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_822 = 7'h36 == predictor_idx_6[6:0] ? predictor_54 : _GEN_821; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_823 = 7'h37 == predictor_idx_6[6:0] ? predictor_55 : _GEN_822; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_824 = 7'h38 == predictor_idx_6[6:0] ? predictor_56 : _GEN_823; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_825 = 7'h39 == predictor_idx_6[6:0] ? predictor_57 : _GEN_824; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_826 = 7'h3a == predictor_idx_6[6:0] ? predictor_58 : _GEN_825; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_827 = 7'h3b == predictor_idx_6[6:0] ? predictor_59 : _GEN_826; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_828 = 7'h3c == predictor_idx_6[6:0] ? predictor_60 : _GEN_827; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_829 = 7'h3d == predictor_idx_6[6:0] ? predictor_61 : _GEN_828; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_830 = 7'h3e == predictor_idx_6[6:0] ? predictor_62 : _GEN_829; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_831 = 7'h3f == predictor_idx_6[6:0] ? predictor_63 : _GEN_830; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_832 = 7'h40 == predictor_idx_6[6:0] ? predictor_64 : _GEN_831; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_833 = 7'h41 == predictor_idx_6[6:0] ? predictor_65 : _GEN_832; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_834 = 7'h42 == predictor_idx_6[6:0] ? predictor_66 : _GEN_833; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_835 = 7'h43 == predictor_idx_6[6:0] ? predictor_67 : _GEN_834; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_836 = 7'h44 == predictor_idx_6[6:0] ? predictor_68 : _GEN_835; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_837 = 7'h45 == predictor_idx_6[6:0] ? predictor_69 : _GEN_836; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_838 = 7'h46 == predictor_idx_6[6:0] ? predictor_70 : _GEN_837; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_839 = 7'h47 == predictor_idx_6[6:0] ? predictor_71 : _GEN_838; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_840 = 7'h48 == predictor_idx_6[6:0] ? predictor_72 : _GEN_839; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_841 = 7'h49 == predictor_idx_6[6:0] ? predictor_73 : _GEN_840; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_842 = 7'h4a == predictor_idx_6[6:0] ? predictor_74 : _GEN_841; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_843 = 7'h4b == predictor_idx_6[6:0] ? predictor_75 : _GEN_842; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_844 = 7'h4c == predictor_idx_6[6:0] ? predictor_76 : _GEN_843; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_845 = 7'h4d == predictor_idx_6[6:0] ? predictor_77 : _GEN_844; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_846 = 7'h4e == predictor_idx_6[6:0] ? predictor_78 : _GEN_845; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_847 = 7'h4f == predictor_idx_6[6:0] ? predictor_79 : _GEN_846; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_848 = 7'h50 == predictor_idx_6[6:0] ? predictor_80 : _GEN_847; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_849 = 7'h51 == predictor_idx_6[6:0] ? predictor_81 : _GEN_848; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_850 = 7'h52 == predictor_idx_6[6:0] ? predictor_82 : _GEN_849; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_851 = 7'h53 == predictor_idx_6[6:0] ? predictor_83 : _GEN_850; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_852 = 7'h54 == predictor_idx_6[6:0] ? predictor_84 : _GEN_851; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_853 = 7'h55 == predictor_idx_6[6:0] ? predictor_85 : _GEN_852; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_854 = 7'h56 == predictor_idx_6[6:0] ? predictor_86 : _GEN_853; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_855 = 7'h57 == predictor_idx_6[6:0] ? predictor_87 : _GEN_854; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_856 = 7'h58 == predictor_idx_6[6:0] ? predictor_88 : _GEN_855; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_857 = 7'h59 == predictor_idx_6[6:0] ? predictor_89 : _GEN_856; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_858 = 7'h5a == predictor_idx_6[6:0] ? predictor_90 : _GEN_857; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_859 = 7'h5b == predictor_idx_6[6:0] ? predictor_91 : _GEN_858; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_860 = 7'h5c == predictor_idx_6[6:0] ? predictor_92 : _GEN_859; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_861 = 7'h5d == predictor_idx_6[6:0] ? predictor_93 : _GEN_860; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_862 = 7'h5e == predictor_idx_6[6:0] ? predictor_94 : _GEN_861; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_863 = 7'h5f == predictor_idx_6[6:0] ? predictor_95 : _GEN_862; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_864 = 7'h60 == predictor_idx_6[6:0] ? predictor_96 : _GEN_863; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_865 = 7'h61 == predictor_idx_6[6:0] ? predictor_97 : _GEN_864; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_866 = 7'h62 == predictor_idx_6[6:0] ? predictor_98 : _GEN_865; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_867 = 7'h63 == predictor_idx_6[6:0] ? predictor_99 : _GEN_866; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_868 = 7'h64 == predictor_idx_6[6:0] ? predictor_100 : _GEN_867; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_869 = 7'h65 == predictor_idx_6[6:0] ? predictor_101 : _GEN_868; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_870 = 7'h66 == predictor_idx_6[6:0] ? predictor_102 : _GEN_869; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_871 = 7'h67 == predictor_idx_6[6:0] ? predictor_103 : _GEN_870; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_872 = 7'h68 == predictor_idx_6[6:0] ? predictor_104 : _GEN_871; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_873 = 7'h69 == predictor_idx_6[6:0] ? predictor_105 : _GEN_872; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_874 = 7'h6a == predictor_idx_6[6:0] ? predictor_106 : _GEN_873; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_875 = 7'h6b == predictor_idx_6[6:0] ? predictor_107 : _GEN_874; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_876 = 7'h6c == predictor_idx_6[6:0] ? predictor_108 : _GEN_875; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_877 = 7'h6d == predictor_idx_6[6:0] ? predictor_109 : _GEN_876; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_878 = 7'h6e == predictor_idx_6[6:0] ? predictor_110 : _GEN_877; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_879 = 7'h6f == predictor_idx_6[6:0] ? predictor_111 : _GEN_878; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_880 = 7'h70 == predictor_idx_6[6:0] ? predictor_112 : _GEN_879; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_881 = 7'h71 == predictor_idx_6[6:0] ? predictor_113 : _GEN_880; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_882 = 7'h72 == predictor_idx_6[6:0] ? predictor_114 : _GEN_881; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_883 = 7'h73 == predictor_idx_6[6:0] ? predictor_115 : _GEN_882; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_884 = 7'h74 == predictor_idx_6[6:0] ? predictor_116 : _GEN_883; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_885 = 7'h75 == predictor_idx_6[6:0] ? predictor_117 : _GEN_884; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_886 = 7'h76 == predictor_idx_6[6:0] ? predictor_118 : _GEN_885; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_887 = 7'h77 == predictor_idx_6[6:0] ? predictor_119 : _GEN_886; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_888 = 7'h78 == predictor_idx_6[6:0] ? predictor_120 : _GEN_887; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_889 = 7'h79 == predictor_idx_6[6:0] ? predictor_121 : _GEN_888; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_890 = 7'h7a == predictor_idx_6[6:0] ? predictor_122 : _GEN_889; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_891 = 7'h7b == predictor_idx_6[6:0] ? predictor_123 : _GEN_890; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_892 = 7'h7c == predictor_idx_6[6:0] ? predictor_124 : _GEN_891; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_893 = 7'h7d == predictor_idx_6[6:0] ? predictor_125 : _GEN_892; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_894 = 7'h7e == predictor_idx_6[6:0] ? predictor_126 : _GEN_893; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_895 = 7'h7f == predictor_idx_6[6:0] ? predictor_127 : _GEN_894; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire  predict_mask_6 = _GEN_895[1]; // @[Bpu.scala 96:62]
  wire [1:0] _GEN_897 = 7'h1 == predictor_idx_7[6:0] ? predictor_1 : predictor_0; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_898 = 7'h2 == predictor_idx_7[6:0] ? predictor_2 : _GEN_897; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_899 = 7'h3 == predictor_idx_7[6:0] ? predictor_3 : _GEN_898; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_900 = 7'h4 == predictor_idx_7[6:0] ? predictor_4 : _GEN_899; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_901 = 7'h5 == predictor_idx_7[6:0] ? predictor_5 : _GEN_900; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_902 = 7'h6 == predictor_idx_7[6:0] ? predictor_6 : _GEN_901; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_903 = 7'h7 == predictor_idx_7[6:0] ? predictor_7 : _GEN_902; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_904 = 7'h8 == predictor_idx_7[6:0] ? predictor_8 : _GEN_903; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_905 = 7'h9 == predictor_idx_7[6:0] ? predictor_9 : _GEN_904; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_906 = 7'ha == predictor_idx_7[6:0] ? predictor_10 : _GEN_905; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_907 = 7'hb == predictor_idx_7[6:0] ? predictor_11 : _GEN_906; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_908 = 7'hc == predictor_idx_7[6:0] ? predictor_12 : _GEN_907; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_909 = 7'hd == predictor_idx_7[6:0] ? predictor_13 : _GEN_908; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_910 = 7'he == predictor_idx_7[6:0] ? predictor_14 : _GEN_909; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_911 = 7'hf == predictor_idx_7[6:0] ? predictor_15 : _GEN_910; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_912 = 7'h10 == predictor_idx_7[6:0] ? predictor_16 : _GEN_911; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_913 = 7'h11 == predictor_idx_7[6:0] ? predictor_17 : _GEN_912; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_914 = 7'h12 == predictor_idx_7[6:0] ? predictor_18 : _GEN_913; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_915 = 7'h13 == predictor_idx_7[6:0] ? predictor_19 : _GEN_914; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_916 = 7'h14 == predictor_idx_7[6:0] ? predictor_20 : _GEN_915; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_917 = 7'h15 == predictor_idx_7[6:0] ? predictor_21 : _GEN_916; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_918 = 7'h16 == predictor_idx_7[6:0] ? predictor_22 : _GEN_917; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_919 = 7'h17 == predictor_idx_7[6:0] ? predictor_23 : _GEN_918; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_920 = 7'h18 == predictor_idx_7[6:0] ? predictor_24 : _GEN_919; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_921 = 7'h19 == predictor_idx_7[6:0] ? predictor_25 : _GEN_920; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_922 = 7'h1a == predictor_idx_7[6:0] ? predictor_26 : _GEN_921; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_923 = 7'h1b == predictor_idx_7[6:0] ? predictor_27 : _GEN_922; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_924 = 7'h1c == predictor_idx_7[6:0] ? predictor_28 : _GEN_923; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_925 = 7'h1d == predictor_idx_7[6:0] ? predictor_29 : _GEN_924; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_926 = 7'h1e == predictor_idx_7[6:0] ? predictor_30 : _GEN_925; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_927 = 7'h1f == predictor_idx_7[6:0] ? predictor_31 : _GEN_926; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_928 = 7'h20 == predictor_idx_7[6:0] ? predictor_32 : _GEN_927; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_929 = 7'h21 == predictor_idx_7[6:0] ? predictor_33 : _GEN_928; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_930 = 7'h22 == predictor_idx_7[6:0] ? predictor_34 : _GEN_929; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_931 = 7'h23 == predictor_idx_7[6:0] ? predictor_35 : _GEN_930; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_932 = 7'h24 == predictor_idx_7[6:0] ? predictor_36 : _GEN_931; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_933 = 7'h25 == predictor_idx_7[6:0] ? predictor_37 : _GEN_932; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_934 = 7'h26 == predictor_idx_7[6:0] ? predictor_38 : _GEN_933; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_935 = 7'h27 == predictor_idx_7[6:0] ? predictor_39 : _GEN_934; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_936 = 7'h28 == predictor_idx_7[6:0] ? predictor_40 : _GEN_935; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_937 = 7'h29 == predictor_idx_7[6:0] ? predictor_41 : _GEN_936; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_938 = 7'h2a == predictor_idx_7[6:0] ? predictor_42 : _GEN_937; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_939 = 7'h2b == predictor_idx_7[6:0] ? predictor_43 : _GEN_938; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_940 = 7'h2c == predictor_idx_7[6:0] ? predictor_44 : _GEN_939; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_941 = 7'h2d == predictor_idx_7[6:0] ? predictor_45 : _GEN_940; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_942 = 7'h2e == predictor_idx_7[6:0] ? predictor_46 : _GEN_941; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_943 = 7'h2f == predictor_idx_7[6:0] ? predictor_47 : _GEN_942; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_944 = 7'h30 == predictor_idx_7[6:0] ? predictor_48 : _GEN_943; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_945 = 7'h31 == predictor_idx_7[6:0] ? predictor_49 : _GEN_944; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_946 = 7'h32 == predictor_idx_7[6:0] ? predictor_50 : _GEN_945; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_947 = 7'h33 == predictor_idx_7[6:0] ? predictor_51 : _GEN_946; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_948 = 7'h34 == predictor_idx_7[6:0] ? predictor_52 : _GEN_947; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_949 = 7'h35 == predictor_idx_7[6:0] ? predictor_53 : _GEN_948; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_950 = 7'h36 == predictor_idx_7[6:0] ? predictor_54 : _GEN_949; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_951 = 7'h37 == predictor_idx_7[6:0] ? predictor_55 : _GEN_950; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_952 = 7'h38 == predictor_idx_7[6:0] ? predictor_56 : _GEN_951; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_953 = 7'h39 == predictor_idx_7[6:0] ? predictor_57 : _GEN_952; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_954 = 7'h3a == predictor_idx_7[6:0] ? predictor_58 : _GEN_953; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_955 = 7'h3b == predictor_idx_7[6:0] ? predictor_59 : _GEN_954; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_956 = 7'h3c == predictor_idx_7[6:0] ? predictor_60 : _GEN_955; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_957 = 7'h3d == predictor_idx_7[6:0] ? predictor_61 : _GEN_956; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_958 = 7'h3e == predictor_idx_7[6:0] ? predictor_62 : _GEN_957; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_959 = 7'h3f == predictor_idx_7[6:0] ? predictor_63 : _GEN_958; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_960 = 7'h40 == predictor_idx_7[6:0] ? predictor_64 : _GEN_959; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_961 = 7'h41 == predictor_idx_7[6:0] ? predictor_65 : _GEN_960; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_962 = 7'h42 == predictor_idx_7[6:0] ? predictor_66 : _GEN_961; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_963 = 7'h43 == predictor_idx_7[6:0] ? predictor_67 : _GEN_962; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_964 = 7'h44 == predictor_idx_7[6:0] ? predictor_68 : _GEN_963; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_965 = 7'h45 == predictor_idx_7[6:0] ? predictor_69 : _GEN_964; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_966 = 7'h46 == predictor_idx_7[6:0] ? predictor_70 : _GEN_965; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_967 = 7'h47 == predictor_idx_7[6:0] ? predictor_71 : _GEN_966; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_968 = 7'h48 == predictor_idx_7[6:0] ? predictor_72 : _GEN_967; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_969 = 7'h49 == predictor_idx_7[6:0] ? predictor_73 : _GEN_968; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_970 = 7'h4a == predictor_idx_7[6:0] ? predictor_74 : _GEN_969; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_971 = 7'h4b == predictor_idx_7[6:0] ? predictor_75 : _GEN_970; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_972 = 7'h4c == predictor_idx_7[6:0] ? predictor_76 : _GEN_971; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_973 = 7'h4d == predictor_idx_7[6:0] ? predictor_77 : _GEN_972; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_974 = 7'h4e == predictor_idx_7[6:0] ? predictor_78 : _GEN_973; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_975 = 7'h4f == predictor_idx_7[6:0] ? predictor_79 : _GEN_974; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_976 = 7'h50 == predictor_idx_7[6:0] ? predictor_80 : _GEN_975; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_977 = 7'h51 == predictor_idx_7[6:0] ? predictor_81 : _GEN_976; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_978 = 7'h52 == predictor_idx_7[6:0] ? predictor_82 : _GEN_977; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_979 = 7'h53 == predictor_idx_7[6:0] ? predictor_83 : _GEN_978; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_980 = 7'h54 == predictor_idx_7[6:0] ? predictor_84 : _GEN_979; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_981 = 7'h55 == predictor_idx_7[6:0] ? predictor_85 : _GEN_980; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_982 = 7'h56 == predictor_idx_7[6:0] ? predictor_86 : _GEN_981; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_983 = 7'h57 == predictor_idx_7[6:0] ? predictor_87 : _GEN_982; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_984 = 7'h58 == predictor_idx_7[6:0] ? predictor_88 : _GEN_983; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_985 = 7'h59 == predictor_idx_7[6:0] ? predictor_89 : _GEN_984; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_986 = 7'h5a == predictor_idx_7[6:0] ? predictor_90 : _GEN_985; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_987 = 7'h5b == predictor_idx_7[6:0] ? predictor_91 : _GEN_986; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_988 = 7'h5c == predictor_idx_7[6:0] ? predictor_92 : _GEN_987; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_989 = 7'h5d == predictor_idx_7[6:0] ? predictor_93 : _GEN_988; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_990 = 7'h5e == predictor_idx_7[6:0] ? predictor_94 : _GEN_989; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_991 = 7'h5f == predictor_idx_7[6:0] ? predictor_95 : _GEN_990; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_992 = 7'h60 == predictor_idx_7[6:0] ? predictor_96 : _GEN_991; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_993 = 7'h61 == predictor_idx_7[6:0] ? predictor_97 : _GEN_992; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_994 = 7'h62 == predictor_idx_7[6:0] ? predictor_98 : _GEN_993; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_995 = 7'h63 == predictor_idx_7[6:0] ? predictor_99 : _GEN_994; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_996 = 7'h64 == predictor_idx_7[6:0] ? predictor_100 : _GEN_995; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_997 = 7'h65 == predictor_idx_7[6:0] ? predictor_101 : _GEN_996; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_998 = 7'h66 == predictor_idx_7[6:0] ? predictor_102 : _GEN_997; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_999 = 7'h67 == predictor_idx_7[6:0] ? predictor_103 : _GEN_998; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_1000 = 7'h68 == predictor_idx_7[6:0] ? predictor_104 : _GEN_999; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_1001 = 7'h69 == predictor_idx_7[6:0] ? predictor_105 : _GEN_1000; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_1002 = 7'h6a == predictor_idx_7[6:0] ? predictor_106 : _GEN_1001; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_1003 = 7'h6b == predictor_idx_7[6:0] ? predictor_107 : _GEN_1002; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_1004 = 7'h6c == predictor_idx_7[6:0] ? predictor_108 : _GEN_1003; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_1005 = 7'h6d == predictor_idx_7[6:0] ? predictor_109 : _GEN_1004; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_1006 = 7'h6e == predictor_idx_7[6:0] ? predictor_110 : _GEN_1005; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_1007 = 7'h6f == predictor_idx_7[6:0] ? predictor_111 : _GEN_1006; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_1008 = 7'h70 == predictor_idx_7[6:0] ? predictor_112 : _GEN_1007; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_1009 = 7'h71 == predictor_idx_7[6:0] ? predictor_113 : _GEN_1008; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_1010 = 7'h72 == predictor_idx_7[6:0] ? predictor_114 : _GEN_1009; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_1011 = 7'h73 == predictor_idx_7[6:0] ? predictor_115 : _GEN_1010; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_1012 = 7'h74 == predictor_idx_7[6:0] ? predictor_116 : _GEN_1011; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_1013 = 7'h75 == predictor_idx_7[6:0] ? predictor_117 : _GEN_1012; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_1014 = 7'h76 == predictor_idx_7[6:0] ? predictor_118 : _GEN_1013; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_1015 = 7'h77 == predictor_idx_7[6:0] ? predictor_119 : _GEN_1014; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_1016 = 7'h78 == predictor_idx_7[6:0] ? predictor_120 : _GEN_1015; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_1017 = 7'h79 == predictor_idx_7[6:0] ? predictor_121 : _GEN_1016; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_1018 = 7'h7a == predictor_idx_7[6:0] ? predictor_122 : _GEN_1017; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_1019 = 7'h7b == predictor_idx_7[6:0] ? predictor_123 : _GEN_1018; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_1020 = 7'h7c == predictor_idx_7[6:0] ? predictor_124 : _GEN_1019; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_1021 = 7'h7d == predictor_idx_7[6:0] ? predictor_125 : _GEN_1020; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_1022 = 7'h7e == predictor_idx_7[6:0] ? predictor_126 : _GEN_1021; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire [1:0] _GEN_1023 = 7'h7f == predictor_idx_7[6:0] ? predictor_127 : _GEN_1022; // @[Bpu.scala 96:62 Bpu.scala 96:62]
  wire  predict_mask_7 = _GEN_1023[1]; // @[Bpu.scala 96:62]
  wire  predict_branch_0 = need_predict_0 & predict_mask_0; // @[Bpu.scala 98:69]
  wire  predict_branch_1 = need_predict_1 & predict_mask_1; // @[Bpu.scala 98:69]
  wire  predict_branch_2 = need_predict_2 & predict_mask_2; // @[Bpu.scala 98:69]
  wire  predict_branch_3 = need_predict_3 & predict_mask_3; // @[Bpu.scala 98:69]
  wire  predict_branch_4 = need_predict_4 & predict_mask_4; // @[Bpu.scala 98:69]
  wire  predict_branch_5 = need_predict_5 & predict_mask_5; // @[Bpu.scala 98:69]
  wire  predict_branch_6 = need_predict_6 & predict_mask_6; // @[Bpu.scala 98:69]
  wire  predict_branch_7 = need_predict_7 & predict_mask_7; // @[Bpu.scala 98:69]
  wire [3:0] is_taken_lo = {predict_branch_3,predict_branch_2,predict_branch_1,predict_branch_0}; // @[Bpu.scala 100:48]
  wire [3:0] is_taken_hi = {predict_branch_7,predict_branch_6,predict_branch_5,predict_branch_4}; // @[Bpu.scala 100:48]
  wire [7:0] _is_taken_T = {predict_branch_7,predict_branch_6,predict_branch_5,predict_branch_4,predict_branch_3,
    predict_branch_2,predict_branch_1,predict_branch_0}; // @[Bpu.scala 100:48]
  wire  is_taken = |_is_taken_T; // @[Bpu.scala 100:54]
  wire [7:0] _inst_mask_enc_T = predict_branch_7 ? 8'h80 : 8'h0; // @[Mux.scala 47:69]
  wire [7:0] _inst_mask_enc_T_1 = predict_branch_6 ? 8'h40 : _inst_mask_enc_T; // @[Mux.scala 47:69]
  wire [7:0] _inst_mask_enc_T_2 = predict_branch_5 ? 8'h20 : _inst_mask_enc_T_1; // @[Mux.scala 47:69]
  wire [7:0] _inst_mask_enc_T_3 = predict_branch_4 ? 8'h10 : _inst_mask_enc_T_2; // @[Mux.scala 47:69]
  wire [7:0] _inst_mask_enc_T_4 = predict_branch_3 ? 8'h8 : _inst_mask_enc_T_3; // @[Mux.scala 47:69]
  wire [7:0] _inst_mask_enc_T_5 = predict_branch_2 ? 8'h4 : _inst_mask_enc_T_4; // @[Mux.scala 47:69]
  wire [7:0] _inst_mask_enc_T_6 = predict_branch_1 ? 8'h2 : _inst_mask_enc_T_5; // @[Mux.scala 47:69]
  wire [7:0] inst_mask_enc = predict_branch_0 ? 8'h1 : _inst_mask_enc_T_6; // @[Mux.scala 47:69]
  wire  inst_mask_0 = inst_mask_enc[0]; // @[OneHot.scala 83:30]
  wire  inst_mask_1 = inst_mask_enc[1]; // @[OneHot.scala 83:30]
  wire  inst_mask_2 = inst_mask_enc[2]; // @[OneHot.scala 83:30]
  wire  inst_mask_3 = inst_mask_enc[3]; // @[OneHot.scala 83:30]
  wire  inst_mask_4 = inst_mask_enc[4]; // @[OneHot.scala 83:30]
  wire  inst_mask_5 = inst_mask_enc[5]; // @[OneHot.scala 83:30]
  wire  inst_mask_6 = inst_mask_enc[6]; // @[OneHot.scala 83:30]
  wire  inst_mask_7 = inst_mask_enc[7]; // @[OneHot.scala 83:30]
  wire [7:0] _inst_idx_T = {inst_mask_7,inst_mask_6,inst_mask_5,inst_mask_4,inst_mask_3,inst_mask_2,inst_mask_1,
    inst_mask_0}; // @[Cat.scala 30:58]
  wire [3:0] inst_idx_hi_1 = _inst_idx_T[7:4]; // @[OneHot.scala 30:18]
  wire [3:0] inst_idx_lo_1 = _inst_idx_T[3:0]; // @[OneHot.scala 31:18]
  wire  inst_idx_hi_2 = |inst_idx_hi_1; // @[OneHot.scala 32:14]
  wire [3:0] _inst_idx_T_1 = inst_idx_hi_1 | inst_idx_lo_1; // @[OneHot.scala 32:28]
  wire [1:0] inst_idx_hi_3 = _inst_idx_T_1[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] inst_idx_lo_2 = _inst_idx_T_1[1:0]; // @[OneHot.scala 31:18]
  wire  inst_idx_hi_4 = |inst_idx_hi_3; // @[OneHot.scala 32:14]
  wire [1:0] _inst_idx_T_2 = inst_idx_hi_3 | inst_idx_lo_2; // @[OneHot.scala 32:28]
  wire  inst_idx_lo_3 = _inst_idx_T_2[1]; // @[CircuitMath.scala 30:8]
  wire [2:0] inst_idx = {inst_idx_hi_2,inst_idx_hi_4,inst_idx_lo_3}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_1025 = 3'h1 == inst_idx ? io_inst_packet_i_bits_data_1 : io_inst_packet_i_bits_data_0; // @[Bpu.scala 108:32 Bpu.scala 108:32]
  wire [31:0] _GEN_1026 = 3'h2 == inst_idx ? io_inst_packet_i_bits_data_2 : _GEN_1025; // @[Bpu.scala 108:32 Bpu.scala 108:32]
  wire [31:0] _GEN_1027 = 3'h3 == inst_idx ? io_inst_packet_i_bits_data_3 : _GEN_1026; // @[Bpu.scala 108:32 Bpu.scala 108:32]
  wire [31:0] _GEN_1028 = 3'h4 == inst_idx ? io_inst_packet_i_bits_data_4 : _GEN_1027; // @[Bpu.scala 108:32 Bpu.scala 108:32]
  wire [31:0] _GEN_1029 = 3'h5 == inst_idx ? io_inst_packet_i_bits_data_5 : _GEN_1028; // @[Bpu.scala 108:32 Bpu.scala 108:32]
  wire [31:0] _GEN_1030 = 3'h6 == inst_idx ? io_inst_packet_i_bits_data_6 : _GEN_1029; // @[Bpu.scala 108:32 Bpu.scala 108:32]
  wire [31:0] _GEN_1031 = 3'h7 == inst_idx ? io_inst_packet_i_bits_data_7 : _GEN_1030; // @[Bpu.scala 108:32 Bpu.scala 108:32]
  wire [13:0] b_imm_hi_hi = _GEN_1031[15] ? 14'h3fff : 14'h0; // @[Bitwise.scala 72:12]
  wire [15:0] b_imm_hi_lo = _GEN_1031[15:0]; // @[Bpu.scala 108:43]
  wire [31:0] _predict_addr_T = {b_imm_hi_hi,b_imm_hi_lo,2'h0}; // @[Bpu.scala 110:35]
  wire [26:0] predict_addr_hi_hi = io_inst_packet_i_bits_addr[31:5]; // @[Bpu.scala 110:70]
  wire [31:0] _predict_addr_T_2 = {predict_addr_hi_hi,inst_idx_hi_2,inst_idx_hi_4,inst_idx_lo_3,2'h0}; // @[Bpu.scala 110:123]
  wire [31:0] _predict_addr_T_5 = $signed(_predict_addr_T) + $signed(_predict_addr_T_2); // @[Bpu.scala 110:38]
  wire [2:0] delay_inst_idx = inst_idx + 3'h1; // @[Bpu.scala 115:33]
  wire  take_delay = inst_idx == 3'h7 & is_taken; // @[Bpu.scala 117:53]
  wire  _GEN_1032 = 3'h0 == delay_inst_idx | (inst_mask_0 | (inst_mask_1 | (inst_mask_2 | (inst_mask_3 | (inst_mask_4 |
    (inst_mask_5 | (inst_mask_6 | (inst_mask_7 | ~is_taken)))))))) & fetched_mask_0; // @[Bpu.scala 122:32 Bpu.scala 122:32 Bpu.scala 119:27]
  wire  _GEN_1033 = 3'h1 == delay_inst_idx | (inst_mask_1 | (inst_mask_2 | (inst_mask_3 | (inst_mask_4 | (inst_mask_5 |
    (inst_mask_6 | (inst_mask_7 | ~is_taken))))))) & fetched_mask_1; // @[Bpu.scala 122:32 Bpu.scala 122:32 Bpu.scala 119:27]
  wire  _GEN_1034 = 3'h2 == delay_inst_idx | (inst_mask_2 | (inst_mask_3 | (inst_mask_4 | (inst_mask_5 | (inst_mask_6 |
    (inst_mask_7 | ~is_taken)))))) & fetched_mask_2; // @[Bpu.scala 122:32 Bpu.scala 122:32 Bpu.scala 119:27]
  wire  _GEN_1035 = 3'h3 == delay_inst_idx | (inst_mask_3 | (inst_mask_4 | (inst_mask_5 | (inst_mask_6 | (inst_mask_7 |
    ~is_taken))))) & fetched_mask_3; // @[Bpu.scala 122:32 Bpu.scala 122:32 Bpu.scala 119:27]
  wire  _GEN_1036 = 3'h4 == delay_inst_idx | (inst_mask_4 | (inst_mask_5 | (inst_mask_6 | (inst_mask_7 | ~is_taken))))
     & fetched_mask_4; // @[Bpu.scala 122:32 Bpu.scala 122:32 Bpu.scala 119:27]
  wire  _GEN_1037 = 3'h5 == delay_inst_idx | (inst_mask_5 | (inst_mask_6 | (inst_mask_7 | ~is_taken))) & fetched_mask_5; // @[Bpu.scala 122:32 Bpu.scala 122:32 Bpu.scala 119:27]
  wire  _GEN_1038 = 3'h6 == delay_inst_idx | (inst_mask_6 | (inst_mask_7 | ~is_taken)) & fetched_mask_6; // @[Bpu.scala 122:32 Bpu.scala 122:32 Bpu.scala 119:27]
  wire  _GEN_1039 = 3'h7 == delay_inst_idx | (inst_mask_7 | ~is_taken) & fetched_mask_7; // @[Bpu.scala 122:32 Bpu.scala 122:32 Bpu.scala 119:27]
  wire [2:0] hi_lo = global_history[3:1]; // @[Bpu.scala 125:148]
  wire [3:0] _hi_T_1 = {is_taken,hi_lo}; // @[Cat.scala 30:58]
  wire [3:0] target_predictor_lo = io_branch_info_i_bits_inst_addr[5:2]; // @[Bpu.scala 126:104]
  wire [7:0] _target_predictor_T = {io_branch_info_i_bits_gh_update,target_predictor_lo}; // @[Cat.scala 30:58]
  wire [1:0] _GEN_1049 = 7'h1 == _target_predictor_T[6:0] ? predictor_1 : predictor_0; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1050 = 7'h2 == _target_predictor_T[6:0] ? predictor_2 : _GEN_1049; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1051 = 7'h3 == _target_predictor_T[6:0] ? predictor_3 : _GEN_1050; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1052 = 7'h4 == _target_predictor_T[6:0] ? predictor_4 : _GEN_1051; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1053 = 7'h5 == _target_predictor_T[6:0] ? predictor_5 : _GEN_1052; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1054 = 7'h6 == _target_predictor_T[6:0] ? predictor_6 : _GEN_1053; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1055 = 7'h7 == _target_predictor_T[6:0] ? predictor_7 : _GEN_1054; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1056 = 7'h8 == _target_predictor_T[6:0] ? predictor_8 : _GEN_1055; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1057 = 7'h9 == _target_predictor_T[6:0] ? predictor_9 : _GEN_1056; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1058 = 7'ha == _target_predictor_T[6:0] ? predictor_10 : _GEN_1057; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1059 = 7'hb == _target_predictor_T[6:0] ? predictor_11 : _GEN_1058; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1060 = 7'hc == _target_predictor_T[6:0] ? predictor_12 : _GEN_1059; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1061 = 7'hd == _target_predictor_T[6:0] ? predictor_13 : _GEN_1060; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1062 = 7'he == _target_predictor_T[6:0] ? predictor_14 : _GEN_1061; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1063 = 7'hf == _target_predictor_T[6:0] ? predictor_15 : _GEN_1062; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1064 = 7'h10 == _target_predictor_T[6:0] ? predictor_16 : _GEN_1063; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1065 = 7'h11 == _target_predictor_T[6:0] ? predictor_17 : _GEN_1064; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1066 = 7'h12 == _target_predictor_T[6:0] ? predictor_18 : _GEN_1065; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1067 = 7'h13 == _target_predictor_T[6:0] ? predictor_19 : _GEN_1066; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1068 = 7'h14 == _target_predictor_T[6:0] ? predictor_20 : _GEN_1067; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1069 = 7'h15 == _target_predictor_T[6:0] ? predictor_21 : _GEN_1068; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1070 = 7'h16 == _target_predictor_T[6:0] ? predictor_22 : _GEN_1069; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1071 = 7'h17 == _target_predictor_T[6:0] ? predictor_23 : _GEN_1070; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1072 = 7'h18 == _target_predictor_T[6:0] ? predictor_24 : _GEN_1071; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1073 = 7'h19 == _target_predictor_T[6:0] ? predictor_25 : _GEN_1072; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1074 = 7'h1a == _target_predictor_T[6:0] ? predictor_26 : _GEN_1073; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1075 = 7'h1b == _target_predictor_T[6:0] ? predictor_27 : _GEN_1074; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1076 = 7'h1c == _target_predictor_T[6:0] ? predictor_28 : _GEN_1075; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1077 = 7'h1d == _target_predictor_T[6:0] ? predictor_29 : _GEN_1076; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1078 = 7'h1e == _target_predictor_T[6:0] ? predictor_30 : _GEN_1077; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1079 = 7'h1f == _target_predictor_T[6:0] ? predictor_31 : _GEN_1078; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1080 = 7'h20 == _target_predictor_T[6:0] ? predictor_32 : _GEN_1079; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1081 = 7'h21 == _target_predictor_T[6:0] ? predictor_33 : _GEN_1080; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1082 = 7'h22 == _target_predictor_T[6:0] ? predictor_34 : _GEN_1081; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1083 = 7'h23 == _target_predictor_T[6:0] ? predictor_35 : _GEN_1082; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1084 = 7'h24 == _target_predictor_T[6:0] ? predictor_36 : _GEN_1083; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1085 = 7'h25 == _target_predictor_T[6:0] ? predictor_37 : _GEN_1084; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1086 = 7'h26 == _target_predictor_T[6:0] ? predictor_38 : _GEN_1085; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1087 = 7'h27 == _target_predictor_T[6:0] ? predictor_39 : _GEN_1086; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1088 = 7'h28 == _target_predictor_T[6:0] ? predictor_40 : _GEN_1087; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1089 = 7'h29 == _target_predictor_T[6:0] ? predictor_41 : _GEN_1088; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1090 = 7'h2a == _target_predictor_T[6:0] ? predictor_42 : _GEN_1089; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1091 = 7'h2b == _target_predictor_T[6:0] ? predictor_43 : _GEN_1090; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1092 = 7'h2c == _target_predictor_T[6:0] ? predictor_44 : _GEN_1091; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1093 = 7'h2d == _target_predictor_T[6:0] ? predictor_45 : _GEN_1092; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1094 = 7'h2e == _target_predictor_T[6:0] ? predictor_46 : _GEN_1093; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1095 = 7'h2f == _target_predictor_T[6:0] ? predictor_47 : _GEN_1094; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1096 = 7'h30 == _target_predictor_T[6:0] ? predictor_48 : _GEN_1095; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1097 = 7'h31 == _target_predictor_T[6:0] ? predictor_49 : _GEN_1096; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1098 = 7'h32 == _target_predictor_T[6:0] ? predictor_50 : _GEN_1097; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1099 = 7'h33 == _target_predictor_T[6:0] ? predictor_51 : _GEN_1098; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1100 = 7'h34 == _target_predictor_T[6:0] ? predictor_52 : _GEN_1099; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1101 = 7'h35 == _target_predictor_T[6:0] ? predictor_53 : _GEN_1100; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1102 = 7'h36 == _target_predictor_T[6:0] ? predictor_54 : _GEN_1101; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1103 = 7'h37 == _target_predictor_T[6:0] ? predictor_55 : _GEN_1102; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1104 = 7'h38 == _target_predictor_T[6:0] ? predictor_56 : _GEN_1103; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1105 = 7'h39 == _target_predictor_T[6:0] ? predictor_57 : _GEN_1104; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1106 = 7'h3a == _target_predictor_T[6:0] ? predictor_58 : _GEN_1105; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1107 = 7'h3b == _target_predictor_T[6:0] ? predictor_59 : _GEN_1106; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1108 = 7'h3c == _target_predictor_T[6:0] ? predictor_60 : _GEN_1107; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1109 = 7'h3d == _target_predictor_T[6:0] ? predictor_61 : _GEN_1108; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1110 = 7'h3e == _target_predictor_T[6:0] ? predictor_62 : _GEN_1109; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1111 = 7'h3f == _target_predictor_T[6:0] ? predictor_63 : _GEN_1110; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1112 = 7'h40 == _target_predictor_T[6:0] ? predictor_64 : _GEN_1111; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1113 = 7'h41 == _target_predictor_T[6:0] ? predictor_65 : _GEN_1112; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1114 = 7'h42 == _target_predictor_T[6:0] ? predictor_66 : _GEN_1113; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1115 = 7'h43 == _target_predictor_T[6:0] ? predictor_67 : _GEN_1114; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1116 = 7'h44 == _target_predictor_T[6:0] ? predictor_68 : _GEN_1115; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1117 = 7'h45 == _target_predictor_T[6:0] ? predictor_69 : _GEN_1116; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1118 = 7'h46 == _target_predictor_T[6:0] ? predictor_70 : _GEN_1117; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1119 = 7'h47 == _target_predictor_T[6:0] ? predictor_71 : _GEN_1118; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1120 = 7'h48 == _target_predictor_T[6:0] ? predictor_72 : _GEN_1119; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1121 = 7'h49 == _target_predictor_T[6:0] ? predictor_73 : _GEN_1120; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1122 = 7'h4a == _target_predictor_T[6:0] ? predictor_74 : _GEN_1121; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1123 = 7'h4b == _target_predictor_T[6:0] ? predictor_75 : _GEN_1122; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1124 = 7'h4c == _target_predictor_T[6:0] ? predictor_76 : _GEN_1123; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1125 = 7'h4d == _target_predictor_T[6:0] ? predictor_77 : _GEN_1124; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1126 = 7'h4e == _target_predictor_T[6:0] ? predictor_78 : _GEN_1125; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1127 = 7'h4f == _target_predictor_T[6:0] ? predictor_79 : _GEN_1126; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1128 = 7'h50 == _target_predictor_T[6:0] ? predictor_80 : _GEN_1127; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1129 = 7'h51 == _target_predictor_T[6:0] ? predictor_81 : _GEN_1128; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1130 = 7'h52 == _target_predictor_T[6:0] ? predictor_82 : _GEN_1129; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1131 = 7'h53 == _target_predictor_T[6:0] ? predictor_83 : _GEN_1130; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1132 = 7'h54 == _target_predictor_T[6:0] ? predictor_84 : _GEN_1131; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1133 = 7'h55 == _target_predictor_T[6:0] ? predictor_85 : _GEN_1132; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1134 = 7'h56 == _target_predictor_T[6:0] ? predictor_86 : _GEN_1133; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1135 = 7'h57 == _target_predictor_T[6:0] ? predictor_87 : _GEN_1134; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1136 = 7'h58 == _target_predictor_T[6:0] ? predictor_88 : _GEN_1135; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1137 = 7'h59 == _target_predictor_T[6:0] ? predictor_89 : _GEN_1136; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1138 = 7'h5a == _target_predictor_T[6:0] ? predictor_90 : _GEN_1137; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1139 = 7'h5b == _target_predictor_T[6:0] ? predictor_91 : _GEN_1138; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1140 = 7'h5c == _target_predictor_T[6:0] ? predictor_92 : _GEN_1139; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1141 = 7'h5d == _target_predictor_T[6:0] ? predictor_93 : _GEN_1140; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1142 = 7'h5e == _target_predictor_T[6:0] ? predictor_94 : _GEN_1141; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1143 = 7'h5f == _target_predictor_T[6:0] ? predictor_95 : _GEN_1142; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1144 = 7'h60 == _target_predictor_T[6:0] ? predictor_96 : _GEN_1143; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1145 = 7'h61 == _target_predictor_T[6:0] ? predictor_97 : _GEN_1144; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1146 = 7'h62 == _target_predictor_T[6:0] ? predictor_98 : _GEN_1145; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1147 = 7'h63 == _target_predictor_T[6:0] ? predictor_99 : _GEN_1146; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1148 = 7'h64 == _target_predictor_T[6:0] ? predictor_100 : _GEN_1147; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1149 = 7'h65 == _target_predictor_T[6:0] ? predictor_101 : _GEN_1148; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1150 = 7'h66 == _target_predictor_T[6:0] ? predictor_102 : _GEN_1149; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1151 = 7'h67 == _target_predictor_T[6:0] ? predictor_103 : _GEN_1150; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1152 = 7'h68 == _target_predictor_T[6:0] ? predictor_104 : _GEN_1151; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1153 = 7'h69 == _target_predictor_T[6:0] ? predictor_105 : _GEN_1152; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1154 = 7'h6a == _target_predictor_T[6:0] ? predictor_106 : _GEN_1153; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1155 = 7'h6b == _target_predictor_T[6:0] ? predictor_107 : _GEN_1154; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1156 = 7'h6c == _target_predictor_T[6:0] ? predictor_108 : _GEN_1155; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1157 = 7'h6d == _target_predictor_T[6:0] ? predictor_109 : _GEN_1156; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1158 = 7'h6e == _target_predictor_T[6:0] ? predictor_110 : _GEN_1157; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1159 = 7'h6f == _target_predictor_T[6:0] ? predictor_111 : _GEN_1158; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1160 = 7'h70 == _target_predictor_T[6:0] ? predictor_112 : _GEN_1159; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1161 = 7'h71 == _target_predictor_T[6:0] ? predictor_113 : _GEN_1160; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1162 = 7'h72 == _target_predictor_T[6:0] ? predictor_114 : _GEN_1161; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1163 = 7'h73 == _target_predictor_T[6:0] ? predictor_115 : _GEN_1162; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1164 = 7'h74 == _target_predictor_T[6:0] ? predictor_116 : _GEN_1163; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1165 = 7'h75 == _target_predictor_T[6:0] ? predictor_117 : _GEN_1164; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1166 = 7'h76 == _target_predictor_T[6:0] ? predictor_118 : _GEN_1165; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1167 = 7'h77 == _target_predictor_T[6:0] ? predictor_119 : _GEN_1166; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1168 = 7'h78 == _target_predictor_T[6:0] ? predictor_120 : _GEN_1167; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1169 = 7'h79 == _target_predictor_T[6:0] ? predictor_121 : _GEN_1168; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1170 = 7'h7a == _target_predictor_T[6:0] ? predictor_122 : _GEN_1169; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1171 = 7'h7b == _target_predictor_T[6:0] ? predictor_123 : _GEN_1170; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1172 = 7'h7c == _target_predictor_T[6:0] ? predictor_124 : _GEN_1171; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1173 = 7'h7d == _target_predictor_T[6:0] ? predictor_125 : _GEN_1172; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1174 = 7'h7e == _target_predictor_T[6:0] ? predictor_126 : _GEN_1173; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire [1:0] _GEN_1175 = 7'h7f == _target_predictor_T[6:0] ? predictor_127 : _GEN_1174; // @[Conditional.scala 37:30 Conditional.scala 37:30]
  wire  _T_3 = 2'h0 == _GEN_1175; // @[Conditional.scala 37:30]
  wire [1:0] _GEN_1176 = 7'h0 == _target_predictor_T[6:0] ? 2'h1 : predictor_0; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1177 = 7'h1 == _target_predictor_T[6:0] ? 2'h1 : predictor_1; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1178 = 7'h2 == _target_predictor_T[6:0] ? 2'h1 : predictor_2; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1179 = 7'h3 == _target_predictor_T[6:0] ? 2'h1 : predictor_3; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1180 = 7'h4 == _target_predictor_T[6:0] ? 2'h1 : predictor_4; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1181 = 7'h5 == _target_predictor_T[6:0] ? 2'h1 : predictor_5; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1182 = 7'h6 == _target_predictor_T[6:0] ? 2'h1 : predictor_6; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1183 = 7'h7 == _target_predictor_T[6:0] ? 2'h1 : predictor_7; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1184 = 7'h8 == _target_predictor_T[6:0] ? 2'h1 : predictor_8; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1185 = 7'h9 == _target_predictor_T[6:0] ? 2'h1 : predictor_9; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1186 = 7'ha == _target_predictor_T[6:0] ? 2'h1 : predictor_10; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1187 = 7'hb == _target_predictor_T[6:0] ? 2'h1 : predictor_11; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1188 = 7'hc == _target_predictor_T[6:0] ? 2'h1 : predictor_12; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1189 = 7'hd == _target_predictor_T[6:0] ? 2'h1 : predictor_13; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1190 = 7'he == _target_predictor_T[6:0] ? 2'h1 : predictor_14; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1191 = 7'hf == _target_predictor_T[6:0] ? 2'h1 : predictor_15; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1192 = 7'h10 == _target_predictor_T[6:0] ? 2'h1 : predictor_16; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1193 = 7'h11 == _target_predictor_T[6:0] ? 2'h1 : predictor_17; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1194 = 7'h12 == _target_predictor_T[6:0] ? 2'h1 : predictor_18; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1195 = 7'h13 == _target_predictor_T[6:0] ? 2'h1 : predictor_19; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1196 = 7'h14 == _target_predictor_T[6:0] ? 2'h1 : predictor_20; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1197 = 7'h15 == _target_predictor_T[6:0] ? 2'h1 : predictor_21; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1198 = 7'h16 == _target_predictor_T[6:0] ? 2'h1 : predictor_22; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1199 = 7'h17 == _target_predictor_T[6:0] ? 2'h1 : predictor_23; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1200 = 7'h18 == _target_predictor_T[6:0] ? 2'h1 : predictor_24; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1201 = 7'h19 == _target_predictor_T[6:0] ? 2'h1 : predictor_25; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1202 = 7'h1a == _target_predictor_T[6:0] ? 2'h1 : predictor_26; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1203 = 7'h1b == _target_predictor_T[6:0] ? 2'h1 : predictor_27; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1204 = 7'h1c == _target_predictor_T[6:0] ? 2'h1 : predictor_28; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1205 = 7'h1d == _target_predictor_T[6:0] ? 2'h1 : predictor_29; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1206 = 7'h1e == _target_predictor_T[6:0] ? 2'h1 : predictor_30; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1207 = 7'h1f == _target_predictor_T[6:0] ? 2'h1 : predictor_31; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1208 = 7'h20 == _target_predictor_T[6:0] ? 2'h1 : predictor_32; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1209 = 7'h21 == _target_predictor_T[6:0] ? 2'h1 : predictor_33; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1210 = 7'h22 == _target_predictor_T[6:0] ? 2'h1 : predictor_34; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1211 = 7'h23 == _target_predictor_T[6:0] ? 2'h1 : predictor_35; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1212 = 7'h24 == _target_predictor_T[6:0] ? 2'h1 : predictor_36; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1213 = 7'h25 == _target_predictor_T[6:0] ? 2'h1 : predictor_37; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1214 = 7'h26 == _target_predictor_T[6:0] ? 2'h1 : predictor_38; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1215 = 7'h27 == _target_predictor_T[6:0] ? 2'h1 : predictor_39; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1216 = 7'h28 == _target_predictor_T[6:0] ? 2'h1 : predictor_40; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1217 = 7'h29 == _target_predictor_T[6:0] ? 2'h1 : predictor_41; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1218 = 7'h2a == _target_predictor_T[6:0] ? 2'h1 : predictor_42; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1219 = 7'h2b == _target_predictor_T[6:0] ? 2'h1 : predictor_43; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1220 = 7'h2c == _target_predictor_T[6:0] ? 2'h1 : predictor_44; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1221 = 7'h2d == _target_predictor_T[6:0] ? 2'h1 : predictor_45; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1222 = 7'h2e == _target_predictor_T[6:0] ? 2'h1 : predictor_46; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1223 = 7'h2f == _target_predictor_T[6:0] ? 2'h1 : predictor_47; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1224 = 7'h30 == _target_predictor_T[6:0] ? 2'h1 : predictor_48; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1225 = 7'h31 == _target_predictor_T[6:0] ? 2'h1 : predictor_49; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1226 = 7'h32 == _target_predictor_T[6:0] ? 2'h1 : predictor_50; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1227 = 7'h33 == _target_predictor_T[6:0] ? 2'h1 : predictor_51; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1228 = 7'h34 == _target_predictor_T[6:0] ? 2'h1 : predictor_52; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1229 = 7'h35 == _target_predictor_T[6:0] ? 2'h1 : predictor_53; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1230 = 7'h36 == _target_predictor_T[6:0] ? 2'h1 : predictor_54; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1231 = 7'h37 == _target_predictor_T[6:0] ? 2'h1 : predictor_55; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1232 = 7'h38 == _target_predictor_T[6:0] ? 2'h1 : predictor_56; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1233 = 7'h39 == _target_predictor_T[6:0] ? 2'h1 : predictor_57; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1234 = 7'h3a == _target_predictor_T[6:0] ? 2'h1 : predictor_58; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1235 = 7'h3b == _target_predictor_T[6:0] ? 2'h1 : predictor_59; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1236 = 7'h3c == _target_predictor_T[6:0] ? 2'h1 : predictor_60; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1237 = 7'h3d == _target_predictor_T[6:0] ? 2'h1 : predictor_61; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1238 = 7'h3e == _target_predictor_T[6:0] ? 2'h1 : predictor_62; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1239 = 7'h3f == _target_predictor_T[6:0] ? 2'h1 : predictor_63; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1240 = 7'h40 == _target_predictor_T[6:0] ? 2'h1 : predictor_64; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1241 = 7'h41 == _target_predictor_T[6:0] ? 2'h1 : predictor_65; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1242 = 7'h42 == _target_predictor_T[6:0] ? 2'h1 : predictor_66; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1243 = 7'h43 == _target_predictor_T[6:0] ? 2'h1 : predictor_67; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1244 = 7'h44 == _target_predictor_T[6:0] ? 2'h1 : predictor_68; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1245 = 7'h45 == _target_predictor_T[6:0] ? 2'h1 : predictor_69; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1246 = 7'h46 == _target_predictor_T[6:0] ? 2'h1 : predictor_70; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1247 = 7'h47 == _target_predictor_T[6:0] ? 2'h1 : predictor_71; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1248 = 7'h48 == _target_predictor_T[6:0] ? 2'h1 : predictor_72; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1249 = 7'h49 == _target_predictor_T[6:0] ? 2'h1 : predictor_73; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1250 = 7'h4a == _target_predictor_T[6:0] ? 2'h1 : predictor_74; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1251 = 7'h4b == _target_predictor_T[6:0] ? 2'h1 : predictor_75; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1252 = 7'h4c == _target_predictor_T[6:0] ? 2'h1 : predictor_76; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1253 = 7'h4d == _target_predictor_T[6:0] ? 2'h1 : predictor_77; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1254 = 7'h4e == _target_predictor_T[6:0] ? 2'h1 : predictor_78; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1255 = 7'h4f == _target_predictor_T[6:0] ? 2'h1 : predictor_79; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1256 = 7'h50 == _target_predictor_T[6:0] ? 2'h1 : predictor_80; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1257 = 7'h51 == _target_predictor_T[6:0] ? 2'h1 : predictor_81; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1258 = 7'h52 == _target_predictor_T[6:0] ? 2'h1 : predictor_82; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1259 = 7'h53 == _target_predictor_T[6:0] ? 2'h1 : predictor_83; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1260 = 7'h54 == _target_predictor_T[6:0] ? 2'h1 : predictor_84; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1261 = 7'h55 == _target_predictor_T[6:0] ? 2'h1 : predictor_85; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1262 = 7'h56 == _target_predictor_T[6:0] ? 2'h1 : predictor_86; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1263 = 7'h57 == _target_predictor_T[6:0] ? 2'h1 : predictor_87; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1264 = 7'h58 == _target_predictor_T[6:0] ? 2'h1 : predictor_88; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1265 = 7'h59 == _target_predictor_T[6:0] ? 2'h1 : predictor_89; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1266 = 7'h5a == _target_predictor_T[6:0] ? 2'h1 : predictor_90; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1267 = 7'h5b == _target_predictor_T[6:0] ? 2'h1 : predictor_91; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1268 = 7'h5c == _target_predictor_T[6:0] ? 2'h1 : predictor_92; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1269 = 7'h5d == _target_predictor_T[6:0] ? 2'h1 : predictor_93; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1270 = 7'h5e == _target_predictor_T[6:0] ? 2'h1 : predictor_94; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1271 = 7'h5f == _target_predictor_T[6:0] ? 2'h1 : predictor_95; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1272 = 7'h60 == _target_predictor_T[6:0] ? 2'h1 : predictor_96; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1273 = 7'h61 == _target_predictor_T[6:0] ? 2'h1 : predictor_97; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1274 = 7'h62 == _target_predictor_T[6:0] ? 2'h1 : predictor_98; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1275 = 7'h63 == _target_predictor_T[6:0] ? 2'h1 : predictor_99; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1276 = 7'h64 == _target_predictor_T[6:0] ? 2'h1 : predictor_100; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1277 = 7'h65 == _target_predictor_T[6:0] ? 2'h1 : predictor_101; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1278 = 7'h66 == _target_predictor_T[6:0] ? 2'h1 : predictor_102; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1279 = 7'h67 == _target_predictor_T[6:0] ? 2'h1 : predictor_103; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1280 = 7'h68 == _target_predictor_T[6:0] ? 2'h1 : predictor_104; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1281 = 7'h69 == _target_predictor_T[6:0] ? 2'h1 : predictor_105; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1282 = 7'h6a == _target_predictor_T[6:0] ? 2'h1 : predictor_106; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1283 = 7'h6b == _target_predictor_T[6:0] ? 2'h1 : predictor_107; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1284 = 7'h6c == _target_predictor_T[6:0] ? 2'h1 : predictor_108; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1285 = 7'h6d == _target_predictor_T[6:0] ? 2'h1 : predictor_109; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1286 = 7'h6e == _target_predictor_T[6:0] ? 2'h1 : predictor_110; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1287 = 7'h6f == _target_predictor_T[6:0] ? 2'h1 : predictor_111; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1288 = 7'h70 == _target_predictor_T[6:0] ? 2'h1 : predictor_112; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1289 = 7'h71 == _target_predictor_T[6:0] ? 2'h1 : predictor_113; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1290 = 7'h72 == _target_predictor_T[6:0] ? 2'h1 : predictor_114; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1291 = 7'h73 == _target_predictor_T[6:0] ? 2'h1 : predictor_115; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1292 = 7'h74 == _target_predictor_T[6:0] ? 2'h1 : predictor_116; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1293 = 7'h75 == _target_predictor_T[6:0] ? 2'h1 : predictor_117; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1294 = 7'h76 == _target_predictor_T[6:0] ? 2'h1 : predictor_118; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1295 = 7'h77 == _target_predictor_T[6:0] ? 2'h1 : predictor_119; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1296 = 7'h78 == _target_predictor_T[6:0] ? 2'h1 : predictor_120; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1297 = 7'h79 == _target_predictor_T[6:0] ? 2'h1 : predictor_121; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1298 = 7'h7a == _target_predictor_T[6:0] ? 2'h1 : predictor_122; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1299 = 7'h7b == _target_predictor_T[6:0] ? 2'h1 : predictor_123; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1300 = 7'h7c == _target_predictor_T[6:0] ? 2'h1 : predictor_124; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1301 = 7'h7d == _target_predictor_T[6:0] ? 2'h1 : predictor_125; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1302 = 7'h7e == _target_predictor_T[6:0] ? 2'h1 : predictor_126; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1303 = 7'h7f == _target_predictor_T[6:0] ? 2'h1 : predictor_127; // @[Bpu.scala 131:28 Bpu.scala 131:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1304 = 7'h0 == _target_predictor_T[6:0] ? 2'h0 : predictor_0; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1305 = 7'h1 == _target_predictor_T[6:0] ? 2'h0 : predictor_1; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1306 = 7'h2 == _target_predictor_T[6:0] ? 2'h0 : predictor_2; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1307 = 7'h3 == _target_predictor_T[6:0] ? 2'h0 : predictor_3; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1308 = 7'h4 == _target_predictor_T[6:0] ? 2'h0 : predictor_4; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1309 = 7'h5 == _target_predictor_T[6:0] ? 2'h0 : predictor_5; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1310 = 7'h6 == _target_predictor_T[6:0] ? 2'h0 : predictor_6; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1311 = 7'h7 == _target_predictor_T[6:0] ? 2'h0 : predictor_7; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1312 = 7'h8 == _target_predictor_T[6:0] ? 2'h0 : predictor_8; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1313 = 7'h9 == _target_predictor_T[6:0] ? 2'h0 : predictor_9; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1314 = 7'ha == _target_predictor_T[6:0] ? 2'h0 : predictor_10; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1315 = 7'hb == _target_predictor_T[6:0] ? 2'h0 : predictor_11; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1316 = 7'hc == _target_predictor_T[6:0] ? 2'h0 : predictor_12; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1317 = 7'hd == _target_predictor_T[6:0] ? 2'h0 : predictor_13; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1318 = 7'he == _target_predictor_T[6:0] ? 2'h0 : predictor_14; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1319 = 7'hf == _target_predictor_T[6:0] ? 2'h0 : predictor_15; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1320 = 7'h10 == _target_predictor_T[6:0] ? 2'h0 : predictor_16; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1321 = 7'h11 == _target_predictor_T[6:0] ? 2'h0 : predictor_17; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1322 = 7'h12 == _target_predictor_T[6:0] ? 2'h0 : predictor_18; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1323 = 7'h13 == _target_predictor_T[6:0] ? 2'h0 : predictor_19; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1324 = 7'h14 == _target_predictor_T[6:0] ? 2'h0 : predictor_20; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1325 = 7'h15 == _target_predictor_T[6:0] ? 2'h0 : predictor_21; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1326 = 7'h16 == _target_predictor_T[6:0] ? 2'h0 : predictor_22; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1327 = 7'h17 == _target_predictor_T[6:0] ? 2'h0 : predictor_23; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1328 = 7'h18 == _target_predictor_T[6:0] ? 2'h0 : predictor_24; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1329 = 7'h19 == _target_predictor_T[6:0] ? 2'h0 : predictor_25; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1330 = 7'h1a == _target_predictor_T[6:0] ? 2'h0 : predictor_26; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1331 = 7'h1b == _target_predictor_T[6:0] ? 2'h0 : predictor_27; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1332 = 7'h1c == _target_predictor_T[6:0] ? 2'h0 : predictor_28; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1333 = 7'h1d == _target_predictor_T[6:0] ? 2'h0 : predictor_29; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1334 = 7'h1e == _target_predictor_T[6:0] ? 2'h0 : predictor_30; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1335 = 7'h1f == _target_predictor_T[6:0] ? 2'h0 : predictor_31; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1336 = 7'h20 == _target_predictor_T[6:0] ? 2'h0 : predictor_32; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1337 = 7'h21 == _target_predictor_T[6:0] ? 2'h0 : predictor_33; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1338 = 7'h22 == _target_predictor_T[6:0] ? 2'h0 : predictor_34; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1339 = 7'h23 == _target_predictor_T[6:0] ? 2'h0 : predictor_35; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1340 = 7'h24 == _target_predictor_T[6:0] ? 2'h0 : predictor_36; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1341 = 7'h25 == _target_predictor_T[6:0] ? 2'h0 : predictor_37; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1342 = 7'h26 == _target_predictor_T[6:0] ? 2'h0 : predictor_38; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1343 = 7'h27 == _target_predictor_T[6:0] ? 2'h0 : predictor_39; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1344 = 7'h28 == _target_predictor_T[6:0] ? 2'h0 : predictor_40; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1345 = 7'h29 == _target_predictor_T[6:0] ? 2'h0 : predictor_41; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1346 = 7'h2a == _target_predictor_T[6:0] ? 2'h0 : predictor_42; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1347 = 7'h2b == _target_predictor_T[6:0] ? 2'h0 : predictor_43; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1348 = 7'h2c == _target_predictor_T[6:0] ? 2'h0 : predictor_44; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1349 = 7'h2d == _target_predictor_T[6:0] ? 2'h0 : predictor_45; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1350 = 7'h2e == _target_predictor_T[6:0] ? 2'h0 : predictor_46; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1351 = 7'h2f == _target_predictor_T[6:0] ? 2'h0 : predictor_47; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1352 = 7'h30 == _target_predictor_T[6:0] ? 2'h0 : predictor_48; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1353 = 7'h31 == _target_predictor_T[6:0] ? 2'h0 : predictor_49; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1354 = 7'h32 == _target_predictor_T[6:0] ? 2'h0 : predictor_50; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1355 = 7'h33 == _target_predictor_T[6:0] ? 2'h0 : predictor_51; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1356 = 7'h34 == _target_predictor_T[6:0] ? 2'h0 : predictor_52; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1357 = 7'h35 == _target_predictor_T[6:0] ? 2'h0 : predictor_53; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1358 = 7'h36 == _target_predictor_T[6:0] ? 2'h0 : predictor_54; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1359 = 7'h37 == _target_predictor_T[6:0] ? 2'h0 : predictor_55; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1360 = 7'h38 == _target_predictor_T[6:0] ? 2'h0 : predictor_56; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1361 = 7'h39 == _target_predictor_T[6:0] ? 2'h0 : predictor_57; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1362 = 7'h3a == _target_predictor_T[6:0] ? 2'h0 : predictor_58; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1363 = 7'h3b == _target_predictor_T[6:0] ? 2'h0 : predictor_59; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1364 = 7'h3c == _target_predictor_T[6:0] ? 2'h0 : predictor_60; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1365 = 7'h3d == _target_predictor_T[6:0] ? 2'h0 : predictor_61; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1366 = 7'h3e == _target_predictor_T[6:0] ? 2'h0 : predictor_62; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1367 = 7'h3f == _target_predictor_T[6:0] ? 2'h0 : predictor_63; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1368 = 7'h40 == _target_predictor_T[6:0] ? 2'h0 : predictor_64; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1369 = 7'h41 == _target_predictor_T[6:0] ? 2'h0 : predictor_65; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1370 = 7'h42 == _target_predictor_T[6:0] ? 2'h0 : predictor_66; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1371 = 7'h43 == _target_predictor_T[6:0] ? 2'h0 : predictor_67; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1372 = 7'h44 == _target_predictor_T[6:0] ? 2'h0 : predictor_68; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1373 = 7'h45 == _target_predictor_T[6:0] ? 2'h0 : predictor_69; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1374 = 7'h46 == _target_predictor_T[6:0] ? 2'h0 : predictor_70; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1375 = 7'h47 == _target_predictor_T[6:0] ? 2'h0 : predictor_71; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1376 = 7'h48 == _target_predictor_T[6:0] ? 2'h0 : predictor_72; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1377 = 7'h49 == _target_predictor_T[6:0] ? 2'h0 : predictor_73; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1378 = 7'h4a == _target_predictor_T[6:0] ? 2'h0 : predictor_74; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1379 = 7'h4b == _target_predictor_T[6:0] ? 2'h0 : predictor_75; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1380 = 7'h4c == _target_predictor_T[6:0] ? 2'h0 : predictor_76; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1381 = 7'h4d == _target_predictor_T[6:0] ? 2'h0 : predictor_77; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1382 = 7'h4e == _target_predictor_T[6:0] ? 2'h0 : predictor_78; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1383 = 7'h4f == _target_predictor_T[6:0] ? 2'h0 : predictor_79; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1384 = 7'h50 == _target_predictor_T[6:0] ? 2'h0 : predictor_80; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1385 = 7'h51 == _target_predictor_T[6:0] ? 2'h0 : predictor_81; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1386 = 7'h52 == _target_predictor_T[6:0] ? 2'h0 : predictor_82; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1387 = 7'h53 == _target_predictor_T[6:0] ? 2'h0 : predictor_83; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1388 = 7'h54 == _target_predictor_T[6:0] ? 2'h0 : predictor_84; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1389 = 7'h55 == _target_predictor_T[6:0] ? 2'h0 : predictor_85; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1390 = 7'h56 == _target_predictor_T[6:0] ? 2'h0 : predictor_86; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1391 = 7'h57 == _target_predictor_T[6:0] ? 2'h0 : predictor_87; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1392 = 7'h58 == _target_predictor_T[6:0] ? 2'h0 : predictor_88; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1393 = 7'h59 == _target_predictor_T[6:0] ? 2'h0 : predictor_89; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1394 = 7'h5a == _target_predictor_T[6:0] ? 2'h0 : predictor_90; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1395 = 7'h5b == _target_predictor_T[6:0] ? 2'h0 : predictor_91; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1396 = 7'h5c == _target_predictor_T[6:0] ? 2'h0 : predictor_92; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1397 = 7'h5d == _target_predictor_T[6:0] ? 2'h0 : predictor_93; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1398 = 7'h5e == _target_predictor_T[6:0] ? 2'h0 : predictor_94; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1399 = 7'h5f == _target_predictor_T[6:0] ? 2'h0 : predictor_95; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1400 = 7'h60 == _target_predictor_T[6:0] ? 2'h0 : predictor_96; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1401 = 7'h61 == _target_predictor_T[6:0] ? 2'h0 : predictor_97; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1402 = 7'h62 == _target_predictor_T[6:0] ? 2'h0 : predictor_98; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1403 = 7'h63 == _target_predictor_T[6:0] ? 2'h0 : predictor_99; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1404 = 7'h64 == _target_predictor_T[6:0] ? 2'h0 : predictor_100; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1405 = 7'h65 == _target_predictor_T[6:0] ? 2'h0 : predictor_101; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1406 = 7'h66 == _target_predictor_T[6:0] ? 2'h0 : predictor_102; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1407 = 7'h67 == _target_predictor_T[6:0] ? 2'h0 : predictor_103; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1408 = 7'h68 == _target_predictor_T[6:0] ? 2'h0 : predictor_104; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1409 = 7'h69 == _target_predictor_T[6:0] ? 2'h0 : predictor_105; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1410 = 7'h6a == _target_predictor_T[6:0] ? 2'h0 : predictor_106; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1411 = 7'h6b == _target_predictor_T[6:0] ? 2'h0 : predictor_107; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1412 = 7'h6c == _target_predictor_T[6:0] ? 2'h0 : predictor_108; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1413 = 7'h6d == _target_predictor_T[6:0] ? 2'h0 : predictor_109; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1414 = 7'h6e == _target_predictor_T[6:0] ? 2'h0 : predictor_110; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1415 = 7'h6f == _target_predictor_T[6:0] ? 2'h0 : predictor_111; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1416 = 7'h70 == _target_predictor_T[6:0] ? 2'h0 : predictor_112; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1417 = 7'h71 == _target_predictor_T[6:0] ? 2'h0 : predictor_113; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1418 = 7'h72 == _target_predictor_T[6:0] ? 2'h0 : predictor_114; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1419 = 7'h73 == _target_predictor_T[6:0] ? 2'h0 : predictor_115; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1420 = 7'h74 == _target_predictor_T[6:0] ? 2'h0 : predictor_116; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1421 = 7'h75 == _target_predictor_T[6:0] ? 2'h0 : predictor_117; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1422 = 7'h76 == _target_predictor_T[6:0] ? 2'h0 : predictor_118; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1423 = 7'h77 == _target_predictor_T[6:0] ? 2'h0 : predictor_119; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1424 = 7'h78 == _target_predictor_T[6:0] ? 2'h0 : predictor_120; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1425 = 7'h79 == _target_predictor_T[6:0] ? 2'h0 : predictor_121; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1426 = 7'h7a == _target_predictor_T[6:0] ? 2'h0 : predictor_122; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1427 = 7'h7b == _target_predictor_T[6:0] ? 2'h0 : predictor_123; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1428 = 7'h7c == _target_predictor_T[6:0] ? 2'h0 : predictor_124; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1429 = 7'h7d == _target_predictor_T[6:0] ? 2'h0 : predictor_125; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1430 = 7'h7e == _target_predictor_T[6:0] ? 2'h0 : predictor_126; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1431 = 7'h7f == _target_predictor_T[6:0] ? 2'h0 : predictor_127; // @[Bpu.scala 133:28 Bpu.scala 133:28 Bpu.scala 74:31]
  wire  _T_4 = 2'h1 == _GEN_1175; // @[Conditional.scala 37:30]
  wire [1:0] _GEN_1560 = 7'h0 == _target_predictor_T[6:0] ? 2'h3 : predictor_0; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1561 = 7'h1 == _target_predictor_T[6:0] ? 2'h3 : predictor_1; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1562 = 7'h2 == _target_predictor_T[6:0] ? 2'h3 : predictor_2; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1563 = 7'h3 == _target_predictor_T[6:0] ? 2'h3 : predictor_3; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1564 = 7'h4 == _target_predictor_T[6:0] ? 2'h3 : predictor_4; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1565 = 7'h5 == _target_predictor_T[6:0] ? 2'h3 : predictor_5; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1566 = 7'h6 == _target_predictor_T[6:0] ? 2'h3 : predictor_6; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1567 = 7'h7 == _target_predictor_T[6:0] ? 2'h3 : predictor_7; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1568 = 7'h8 == _target_predictor_T[6:0] ? 2'h3 : predictor_8; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1569 = 7'h9 == _target_predictor_T[6:0] ? 2'h3 : predictor_9; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1570 = 7'ha == _target_predictor_T[6:0] ? 2'h3 : predictor_10; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1571 = 7'hb == _target_predictor_T[6:0] ? 2'h3 : predictor_11; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1572 = 7'hc == _target_predictor_T[6:0] ? 2'h3 : predictor_12; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1573 = 7'hd == _target_predictor_T[6:0] ? 2'h3 : predictor_13; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1574 = 7'he == _target_predictor_T[6:0] ? 2'h3 : predictor_14; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1575 = 7'hf == _target_predictor_T[6:0] ? 2'h3 : predictor_15; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1576 = 7'h10 == _target_predictor_T[6:0] ? 2'h3 : predictor_16; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1577 = 7'h11 == _target_predictor_T[6:0] ? 2'h3 : predictor_17; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1578 = 7'h12 == _target_predictor_T[6:0] ? 2'h3 : predictor_18; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1579 = 7'h13 == _target_predictor_T[6:0] ? 2'h3 : predictor_19; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1580 = 7'h14 == _target_predictor_T[6:0] ? 2'h3 : predictor_20; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1581 = 7'h15 == _target_predictor_T[6:0] ? 2'h3 : predictor_21; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1582 = 7'h16 == _target_predictor_T[6:0] ? 2'h3 : predictor_22; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1583 = 7'h17 == _target_predictor_T[6:0] ? 2'h3 : predictor_23; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1584 = 7'h18 == _target_predictor_T[6:0] ? 2'h3 : predictor_24; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1585 = 7'h19 == _target_predictor_T[6:0] ? 2'h3 : predictor_25; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1586 = 7'h1a == _target_predictor_T[6:0] ? 2'h3 : predictor_26; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1587 = 7'h1b == _target_predictor_T[6:0] ? 2'h3 : predictor_27; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1588 = 7'h1c == _target_predictor_T[6:0] ? 2'h3 : predictor_28; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1589 = 7'h1d == _target_predictor_T[6:0] ? 2'h3 : predictor_29; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1590 = 7'h1e == _target_predictor_T[6:0] ? 2'h3 : predictor_30; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1591 = 7'h1f == _target_predictor_T[6:0] ? 2'h3 : predictor_31; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1592 = 7'h20 == _target_predictor_T[6:0] ? 2'h3 : predictor_32; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1593 = 7'h21 == _target_predictor_T[6:0] ? 2'h3 : predictor_33; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1594 = 7'h22 == _target_predictor_T[6:0] ? 2'h3 : predictor_34; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1595 = 7'h23 == _target_predictor_T[6:0] ? 2'h3 : predictor_35; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1596 = 7'h24 == _target_predictor_T[6:0] ? 2'h3 : predictor_36; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1597 = 7'h25 == _target_predictor_T[6:0] ? 2'h3 : predictor_37; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1598 = 7'h26 == _target_predictor_T[6:0] ? 2'h3 : predictor_38; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1599 = 7'h27 == _target_predictor_T[6:0] ? 2'h3 : predictor_39; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1600 = 7'h28 == _target_predictor_T[6:0] ? 2'h3 : predictor_40; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1601 = 7'h29 == _target_predictor_T[6:0] ? 2'h3 : predictor_41; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1602 = 7'h2a == _target_predictor_T[6:0] ? 2'h3 : predictor_42; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1603 = 7'h2b == _target_predictor_T[6:0] ? 2'h3 : predictor_43; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1604 = 7'h2c == _target_predictor_T[6:0] ? 2'h3 : predictor_44; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1605 = 7'h2d == _target_predictor_T[6:0] ? 2'h3 : predictor_45; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1606 = 7'h2e == _target_predictor_T[6:0] ? 2'h3 : predictor_46; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1607 = 7'h2f == _target_predictor_T[6:0] ? 2'h3 : predictor_47; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1608 = 7'h30 == _target_predictor_T[6:0] ? 2'h3 : predictor_48; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1609 = 7'h31 == _target_predictor_T[6:0] ? 2'h3 : predictor_49; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1610 = 7'h32 == _target_predictor_T[6:0] ? 2'h3 : predictor_50; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1611 = 7'h33 == _target_predictor_T[6:0] ? 2'h3 : predictor_51; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1612 = 7'h34 == _target_predictor_T[6:0] ? 2'h3 : predictor_52; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1613 = 7'h35 == _target_predictor_T[6:0] ? 2'h3 : predictor_53; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1614 = 7'h36 == _target_predictor_T[6:0] ? 2'h3 : predictor_54; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1615 = 7'h37 == _target_predictor_T[6:0] ? 2'h3 : predictor_55; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1616 = 7'h38 == _target_predictor_T[6:0] ? 2'h3 : predictor_56; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1617 = 7'h39 == _target_predictor_T[6:0] ? 2'h3 : predictor_57; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1618 = 7'h3a == _target_predictor_T[6:0] ? 2'h3 : predictor_58; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1619 = 7'h3b == _target_predictor_T[6:0] ? 2'h3 : predictor_59; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1620 = 7'h3c == _target_predictor_T[6:0] ? 2'h3 : predictor_60; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1621 = 7'h3d == _target_predictor_T[6:0] ? 2'h3 : predictor_61; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1622 = 7'h3e == _target_predictor_T[6:0] ? 2'h3 : predictor_62; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1623 = 7'h3f == _target_predictor_T[6:0] ? 2'h3 : predictor_63; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1624 = 7'h40 == _target_predictor_T[6:0] ? 2'h3 : predictor_64; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1625 = 7'h41 == _target_predictor_T[6:0] ? 2'h3 : predictor_65; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1626 = 7'h42 == _target_predictor_T[6:0] ? 2'h3 : predictor_66; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1627 = 7'h43 == _target_predictor_T[6:0] ? 2'h3 : predictor_67; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1628 = 7'h44 == _target_predictor_T[6:0] ? 2'h3 : predictor_68; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1629 = 7'h45 == _target_predictor_T[6:0] ? 2'h3 : predictor_69; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1630 = 7'h46 == _target_predictor_T[6:0] ? 2'h3 : predictor_70; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1631 = 7'h47 == _target_predictor_T[6:0] ? 2'h3 : predictor_71; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1632 = 7'h48 == _target_predictor_T[6:0] ? 2'h3 : predictor_72; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1633 = 7'h49 == _target_predictor_T[6:0] ? 2'h3 : predictor_73; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1634 = 7'h4a == _target_predictor_T[6:0] ? 2'h3 : predictor_74; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1635 = 7'h4b == _target_predictor_T[6:0] ? 2'h3 : predictor_75; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1636 = 7'h4c == _target_predictor_T[6:0] ? 2'h3 : predictor_76; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1637 = 7'h4d == _target_predictor_T[6:0] ? 2'h3 : predictor_77; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1638 = 7'h4e == _target_predictor_T[6:0] ? 2'h3 : predictor_78; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1639 = 7'h4f == _target_predictor_T[6:0] ? 2'h3 : predictor_79; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1640 = 7'h50 == _target_predictor_T[6:0] ? 2'h3 : predictor_80; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1641 = 7'h51 == _target_predictor_T[6:0] ? 2'h3 : predictor_81; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1642 = 7'h52 == _target_predictor_T[6:0] ? 2'h3 : predictor_82; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1643 = 7'h53 == _target_predictor_T[6:0] ? 2'h3 : predictor_83; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1644 = 7'h54 == _target_predictor_T[6:0] ? 2'h3 : predictor_84; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1645 = 7'h55 == _target_predictor_T[6:0] ? 2'h3 : predictor_85; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1646 = 7'h56 == _target_predictor_T[6:0] ? 2'h3 : predictor_86; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1647 = 7'h57 == _target_predictor_T[6:0] ? 2'h3 : predictor_87; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1648 = 7'h58 == _target_predictor_T[6:0] ? 2'h3 : predictor_88; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1649 = 7'h59 == _target_predictor_T[6:0] ? 2'h3 : predictor_89; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1650 = 7'h5a == _target_predictor_T[6:0] ? 2'h3 : predictor_90; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1651 = 7'h5b == _target_predictor_T[6:0] ? 2'h3 : predictor_91; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1652 = 7'h5c == _target_predictor_T[6:0] ? 2'h3 : predictor_92; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1653 = 7'h5d == _target_predictor_T[6:0] ? 2'h3 : predictor_93; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1654 = 7'h5e == _target_predictor_T[6:0] ? 2'h3 : predictor_94; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1655 = 7'h5f == _target_predictor_T[6:0] ? 2'h3 : predictor_95; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1656 = 7'h60 == _target_predictor_T[6:0] ? 2'h3 : predictor_96; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1657 = 7'h61 == _target_predictor_T[6:0] ? 2'h3 : predictor_97; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1658 = 7'h62 == _target_predictor_T[6:0] ? 2'h3 : predictor_98; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1659 = 7'h63 == _target_predictor_T[6:0] ? 2'h3 : predictor_99; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1660 = 7'h64 == _target_predictor_T[6:0] ? 2'h3 : predictor_100; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1661 = 7'h65 == _target_predictor_T[6:0] ? 2'h3 : predictor_101; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1662 = 7'h66 == _target_predictor_T[6:0] ? 2'h3 : predictor_102; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1663 = 7'h67 == _target_predictor_T[6:0] ? 2'h3 : predictor_103; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1664 = 7'h68 == _target_predictor_T[6:0] ? 2'h3 : predictor_104; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1665 = 7'h69 == _target_predictor_T[6:0] ? 2'h3 : predictor_105; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1666 = 7'h6a == _target_predictor_T[6:0] ? 2'h3 : predictor_106; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1667 = 7'h6b == _target_predictor_T[6:0] ? 2'h3 : predictor_107; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1668 = 7'h6c == _target_predictor_T[6:0] ? 2'h3 : predictor_108; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1669 = 7'h6d == _target_predictor_T[6:0] ? 2'h3 : predictor_109; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1670 = 7'h6e == _target_predictor_T[6:0] ? 2'h3 : predictor_110; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1671 = 7'h6f == _target_predictor_T[6:0] ? 2'h3 : predictor_111; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1672 = 7'h70 == _target_predictor_T[6:0] ? 2'h3 : predictor_112; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1673 = 7'h71 == _target_predictor_T[6:0] ? 2'h3 : predictor_113; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1674 = 7'h72 == _target_predictor_T[6:0] ? 2'h3 : predictor_114; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1675 = 7'h73 == _target_predictor_T[6:0] ? 2'h3 : predictor_115; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1676 = 7'h74 == _target_predictor_T[6:0] ? 2'h3 : predictor_116; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1677 = 7'h75 == _target_predictor_T[6:0] ? 2'h3 : predictor_117; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1678 = 7'h76 == _target_predictor_T[6:0] ? 2'h3 : predictor_118; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1679 = 7'h77 == _target_predictor_T[6:0] ? 2'h3 : predictor_119; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1680 = 7'h78 == _target_predictor_T[6:0] ? 2'h3 : predictor_120; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1681 = 7'h79 == _target_predictor_T[6:0] ? 2'h3 : predictor_121; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1682 = 7'h7a == _target_predictor_T[6:0] ? 2'h3 : predictor_122; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1683 = 7'h7b == _target_predictor_T[6:0] ? 2'h3 : predictor_123; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1684 = 7'h7c == _target_predictor_T[6:0] ? 2'h3 : predictor_124; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1685 = 7'h7d == _target_predictor_T[6:0] ? 2'h3 : predictor_125; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1686 = 7'h7e == _target_predictor_T[6:0] ? 2'h3 : predictor_126; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1687 = 7'h7f == _target_predictor_T[6:0] ? 2'h3 : predictor_127; // @[Bpu.scala 138:28 Bpu.scala 138:28 Bpu.scala 74:31]
  wire [1:0] _GEN_1816 = io_branch_info_i_bits_is_taken ? _GEN_1560 : _GEN_1304; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1817 = io_branch_info_i_bits_is_taken ? _GEN_1561 : _GEN_1305; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1818 = io_branch_info_i_bits_is_taken ? _GEN_1562 : _GEN_1306; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1819 = io_branch_info_i_bits_is_taken ? _GEN_1563 : _GEN_1307; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1820 = io_branch_info_i_bits_is_taken ? _GEN_1564 : _GEN_1308; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1821 = io_branch_info_i_bits_is_taken ? _GEN_1565 : _GEN_1309; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1822 = io_branch_info_i_bits_is_taken ? _GEN_1566 : _GEN_1310; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1823 = io_branch_info_i_bits_is_taken ? _GEN_1567 : _GEN_1311; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1824 = io_branch_info_i_bits_is_taken ? _GEN_1568 : _GEN_1312; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1825 = io_branch_info_i_bits_is_taken ? _GEN_1569 : _GEN_1313; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1826 = io_branch_info_i_bits_is_taken ? _GEN_1570 : _GEN_1314; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1827 = io_branch_info_i_bits_is_taken ? _GEN_1571 : _GEN_1315; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1828 = io_branch_info_i_bits_is_taken ? _GEN_1572 : _GEN_1316; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1829 = io_branch_info_i_bits_is_taken ? _GEN_1573 : _GEN_1317; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1830 = io_branch_info_i_bits_is_taken ? _GEN_1574 : _GEN_1318; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1831 = io_branch_info_i_bits_is_taken ? _GEN_1575 : _GEN_1319; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1832 = io_branch_info_i_bits_is_taken ? _GEN_1576 : _GEN_1320; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1833 = io_branch_info_i_bits_is_taken ? _GEN_1577 : _GEN_1321; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1834 = io_branch_info_i_bits_is_taken ? _GEN_1578 : _GEN_1322; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1835 = io_branch_info_i_bits_is_taken ? _GEN_1579 : _GEN_1323; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1836 = io_branch_info_i_bits_is_taken ? _GEN_1580 : _GEN_1324; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1837 = io_branch_info_i_bits_is_taken ? _GEN_1581 : _GEN_1325; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1838 = io_branch_info_i_bits_is_taken ? _GEN_1582 : _GEN_1326; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1839 = io_branch_info_i_bits_is_taken ? _GEN_1583 : _GEN_1327; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1840 = io_branch_info_i_bits_is_taken ? _GEN_1584 : _GEN_1328; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1841 = io_branch_info_i_bits_is_taken ? _GEN_1585 : _GEN_1329; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1842 = io_branch_info_i_bits_is_taken ? _GEN_1586 : _GEN_1330; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1843 = io_branch_info_i_bits_is_taken ? _GEN_1587 : _GEN_1331; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1844 = io_branch_info_i_bits_is_taken ? _GEN_1588 : _GEN_1332; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1845 = io_branch_info_i_bits_is_taken ? _GEN_1589 : _GEN_1333; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1846 = io_branch_info_i_bits_is_taken ? _GEN_1590 : _GEN_1334; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1847 = io_branch_info_i_bits_is_taken ? _GEN_1591 : _GEN_1335; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1848 = io_branch_info_i_bits_is_taken ? _GEN_1592 : _GEN_1336; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1849 = io_branch_info_i_bits_is_taken ? _GEN_1593 : _GEN_1337; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1850 = io_branch_info_i_bits_is_taken ? _GEN_1594 : _GEN_1338; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1851 = io_branch_info_i_bits_is_taken ? _GEN_1595 : _GEN_1339; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1852 = io_branch_info_i_bits_is_taken ? _GEN_1596 : _GEN_1340; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1853 = io_branch_info_i_bits_is_taken ? _GEN_1597 : _GEN_1341; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1854 = io_branch_info_i_bits_is_taken ? _GEN_1598 : _GEN_1342; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1855 = io_branch_info_i_bits_is_taken ? _GEN_1599 : _GEN_1343; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1856 = io_branch_info_i_bits_is_taken ? _GEN_1600 : _GEN_1344; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1857 = io_branch_info_i_bits_is_taken ? _GEN_1601 : _GEN_1345; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1858 = io_branch_info_i_bits_is_taken ? _GEN_1602 : _GEN_1346; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1859 = io_branch_info_i_bits_is_taken ? _GEN_1603 : _GEN_1347; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1860 = io_branch_info_i_bits_is_taken ? _GEN_1604 : _GEN_1348; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1861 = io_branch_info_i_bits_is_taken ? _GEN_1605 : _GEN_1349; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1862 = io_branch_info_i_bits_is_taken ? _GEN_1606 : _GEN_1350; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1863 = io_branch_info_i_bits_is_taken ? _GEN_1607 : _GEN_1351; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1864 = io_branch_info_i_bits_is_taken ? _GEN_1608 : _GEN_1352; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1865 = io_branch_info_i_bits_is_taken ? _GEN_1609 : _GEN_1353; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1866 = io_branch_info_i_bits_is_taken ? _GEN_1610 : _GEN_1354; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1867 = io_branch_info_i_bits_is_taken ? _GEN_1611 : _GEN_1355; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1868 = io_branch_info_i_bits_is_taken ? _GEN_1612 : _GEN_1356; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1869 = io_branch_info_i_bits_is_taken ? _GEN_1613 : _GEN_1357; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1870 = io_branch_info_i_bits_is_taken ? _GEN_1614 : _GEN_1358; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1871 = io_branch_info_i_bits_is_taken ? _GEN_1615 : _GEN_1359; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1872 = io_branch_info_i_bits_is_taken ? _GEN_1616 : _GEN_1360; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1873 = io_branch_info_i_bits_is_taken ? _GEN_1617 : _GEN_1361; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1874 = io_branch_info_i_bits_is_taken ? _GEN_1618 : _GEN_1362; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1875 = io_branch_info_i_bits_is_taken ? _GEN_1619 : _GEN_1363; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1876 = io_branch_info_i_bits_is_taken ? _GEN_1620 : _GEN_1364; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1877 = io_branch_info_i_bits_is_taken ? _GEN_1621 : _GEN_1365; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1878 = io_branch_info_i_bits_is_taken ? _GEN_1622 : _GEN_1366; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1879 = io_branch_info_i_bits_is_taken ? _GEN_1623 : _GEN_1367; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1880 = io_branch_info_i_bits_is_taken ? _GEN_1624 : _GEN_1368; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1881 = io_branch_info_i_bits_is_taken ? _GEN_1625 : _GEN_1369; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1882 = io_branch_info_i_bits_is_taken ? _GEN_1626 : _GEN_1370; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1883 = io_branch_info_i_bits_is_taken ? _GEN_1627 : _GEN_1371; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1884 = io_branch_info_i_bits_is_taken ? _GEN_1628 : _GEN_1372; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1885 = io_branch_info_i_bits_is_taken ? _GEN_1629 : _GEN_1373; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1886 = io_branch_info_i_bits_is_taken ? _GEN_1630 : _GEN_1374; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1887 = io_branch_info_i_bits_is_taken ? _GEN_1631 : _GEN_1375; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1888 = io_branch_info_i_bits_is_taken ? _GEN_1632 : _GEN_1376; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1889 = io_branch_info_i_bits_is_taken ? _GEN_1633 : _GEN_1377; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1890 = io_branch_info_i_bits_is_taken ? _GEN_1634 : _GEN_1378; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1891 = io_branch_info_i_bits_is_taken ? _GEN_1635 : _GEN_1379; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1892 = io_branch_info_i_bits_is_taken ? _GEN_1636 : _GEN_1380; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1893 = io_branch_info_i_bits_is_taken ? _GEN_1637 : _GEN_1381; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1894 = io_branch_info_i_bits_is_taken ? _GEN_1638 : _GEN_1382; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1895 = io_branch_info_i_bits_is_taken ? _GEN_1639 : _GEN_1383; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1896 = io_branch_info_i_bits_is_taken ? _GEN_1640 : _GEN_1384; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1897 = io_branch_info_i_bits_is_taken ? _GEN_1641 : _GEN_1385; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1898 = io_branch_info_i_bits_is_taken ? _GEN_1642 : _GEN_1386; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1899 = io_branch_info_i_bits_is_taken ? _GEN_1643 : _GEN_1387; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1900 = io_branch_info_i_bits_is_taken ? _GEN_1644 : _GEN_1388; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1901 = io_branch_info_i_bits_is_taken ? _GEN_1645 : _GEN_1389; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1902 = io_branch_info_i_bits_is_taken ? _GEN_1646 : _GEN_1390; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1903 = io_branch_info_i_bits_is_taken ? _GEN_1647 : _GEN_1391; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1904 = io_branch_info_i_bits_is_taken ? _GEN_1648 : _GEN_1392; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1905 = io_branch_info_i_bits_is_taken ? _GEN_1649 : _GEN_1393; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1906 = io_branch_info_i_bits_is_taken ? _GEN_1650 : _GEN_1394; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1907 = io_branch_info_i_bits_is_taken ? _GEN_1651 : _GEN_1395; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1908 = io_branch_info_i_bits_is_taken ? _GEN_1652 : _GEN_1396; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1909 = io_branch_info_i_bits_is_taken ? _GEN_1653 : _GEN_1397; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1910 = io_branch_info_i_bits_is_taken ? _GEN_1654 : _GEN_1398; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1911 = io_branch_info_i_bits_is_taken ? _GEN_1655 : _GEN_1399; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1912 = io_branch_info_i_bits_is_taken ? _GEN_1656 : _GEN_1400; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1913 = io_branch_info_i_bits_is_taken ? _GEN_1657 : _GEN_1401; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1914 = io_branch_info_i_bits_is_taken ? _GEN_1658 : _GEN_1402; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1915 = io_branch_info_i_bits_is_taken ? _GEN_1659 : _GEN_1403; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1916 = io_branch_info_i_bits_is_taken ? _GEN_1660 : _GEN_1404; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1917 = io_branch_info_i_bits_is_taken ? _GEN_1661 : _GEN_1405; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1918 = io_branch_info_i_bits_is_taken ? _GEN_1662 : _GEN_1406; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1919 = io_branch_info_i_bits_is_taken ? _GEN_1663 : _GEN_1407; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1920 = io_branch_info_i_bits_is_taken ? _GEN_1664 : _GEN_1408; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1921 = io_branch_info_i_bits_is_taken ? _GEN_1665 : _GEN_1409; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1922 = io_branch_info_i_bits_is_taken ? _GEN_1666 : _GEN_1410; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1923 = io_branch_info_i_bits_is_taken ? _GEN_1667 : _GEN_1411; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1924 = io_branch_info_i_bits_is_taken ? _GEN_1668 : _GEN_1412; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1925 = io_branch_info_i_bits_is_taken ? _GEN_1669 : _GEN_1413; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1926 = io_branch_info_i_bits_is_taken ? _GEN_1670 : _GEN_1414; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1927 = io_branch_info_i_bits_is_taken ? _GEN_1671 : _GEN_1415; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1928 = io_branch_info_i_bits_is_taken ? _GEN_1672 : _GEN_1416; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1929 = io_branch_info_i_bits_is_taken ? _GEN_1673 : _GEN_1417; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1930 = io_branch_info_i_bits_is_taken ? _GEN_1674 : _GEN_1418; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1931 = io_branch_info_i_bits_is_taken ? _GEN_1675 : _GEN_1419; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1932 = io_branch_info_i_bits_is_taken ? _GEN_1676 : _GEN_1420; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1933 = io_branch_info_i_bits_is_taken ? _GEN_1677 : _GEN_1421; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1934 = io_branch_info_i_bits_is_taken ? _GEN_1678 : _GEN_1422; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1935 = io_branch_info_i_bits_is_taken ? _GEN_1679 : _GEN_1423; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1936 = io_branch_info_i_bits_is_taken ? _GEN_1680 : _GEN_1424; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1937 = io_branch_info_i_bits_is_taken ? _GEN_1681 : _GEN_1425; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1938 = io_branch_info_i_bits_is_taken ? _GEN_1682 : _GEN_1426; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1939 = io_branch_info_i_bits_is_taken ? _GEN_1683 : _GEN_1427; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1940 = io_branch_info_i_bits_is_taken ? _GEN_1684 : _GEN_1428; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1941 = io_branch_info_i_bits_is_taken ? _GEN_1685 : _GEN_1429; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1942 = io_branch_info_i_bits_is_taken ? _GEN_1686 : _GEN_1430; // @[Bpu.scala 137:46]
  wire [1:0] _GEN_1943 = io_branch_info_i_bits_is_taken ? _GEN_1687 : _GEN_1431; // @[Bpu.scala 137:46]
  wire  _T_5 = 2'h2 == _GEN_1175; // @[Conditional.scala 37:30]
  wire  _T_6 = 2'h3 == _GEN_1175; // @[Conditional.scala 37:30]
  wire [1:0] _GEN_2456 = 7'h0 == _target_predictor_T[6:0] ? 2'h2 : predictor_0; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2457 = 7'h1 == _target_predictor_T[6:0] ? 2'h2 : predictor_1; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2458 = 7'h2 == _target_predictor_T[6:0] ? 2'h2 : predictor_2; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2459 = 7'h3 == _target_predictor_T[6:0] ? 2'h2 : predictor_3; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2460 = 7'h4 == _target_predictor_T[6:0] ? 2'h2 : predictor_4; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2461 = 7'h5 == _target_predictor_T[6:0] ? 2'h2 : predictor_5; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2462 = 7'h6 == _target_predictor_T[6:0] ? 2'h2 : predictor_6; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2463 = 7'h7 == _target_predictor_T[6:0] ? 2'h2 : predictor_7; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2464 = 7'h8 == _target_predictor_T[6:0] ? 2'h2 : predictor_8; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2465 = 7'h9 == _target_predictor_T[6:0] ? 2'h2 : predictor_9; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2466 = 7'ha == _target_predictor_T[6:0] ? 2'h2 : predictor_10; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2467 = 7'hb == _target_predictor_T[6:0] ? 2'h2 : predictor_11; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2468 = 7'hc == _target_predictor_T[6:0] ? 2'h2 : predictor_12; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2469 = 7'hd == _target_predictor_T[6:0] ? 2'h2 : predictor_13; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2470 = 7'he == _target_predictor_T[6:0] ? 2'h2 : predictor_14; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2471 = 7'hf == _target_predictor_T[6:0] ? 2'h2 : predictor_15; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2472 = 7'h10 == _target_predictor_T[6:0] ? 2'h2 : predictor_16; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2473 = 7'h11 == _target_predictor_T[6:0] ? 2'h2 : predictor_17; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2474 = 7'h12 == _target_predictor_T[6:0] ? 2'h2 : predictor_18; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2475 = 7'h13 == _target_predictor_T[6:0] ? 2'h2 : predictor_19; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2476 = 7'h14 == _target_predictor_T[6:0] ? 2'h2 : predictor_20; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2477 = 7'h15 == _target_predictor_T[6:0] ? 2'h2 : predictor_21; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2478 = 7'h16 == _target_predictor_T[6:0] ? 2'h2 : predictor_22; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2479 = 7'h17 == _target_predictor_T[6:0] ? 2'h2 : predictor_23; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2480 = 7'h18 == _target_predictor_T[6:0] ? 2'h2 : predictor_24; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2481 = 7'h19 == _target_predictor_T[6:0] ? 2'h2 : predictor_25; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2482 = 7'h1a == _target_predictor_T[6:0] ? 2'h2 : predictor_26; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2483 = 7'h1b == _target_predictor_T[6:0] ? 2'h2 : predictor_27; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2484 = 7'h1c == _target_predictor_T[6:0] ? 2'h2 : predictor_28; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2485 = 7'h1d == _target_predictor_T[6:0] ? 2'h2 : predictor_29; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2486 = 7'h1e == _target_predictor_T[6:0] ? 2'h2 : predictor_30; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2487 = 7'h1f == _target_predictor_T[6:0] ? 2'h2 : predictor_31; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2488 = 7'h20 == _target_predictor_T[6:0] ? 2'h2 : predictor_32; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2489 = 7'h21 == _target_predictor_T[6:0] ? 2'h2 : predictor_33; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2490 = 7'h22 == _target_predictor_T[6:0] ? 2'h2 : predictor_34; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2491 = 7'h23 == _target_predictor_T[6:0] ? 2'h2 : predictor_35; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2492 = 7'h24 == _target_predictor_T[6:0] ? 2'h2 : predictor_36; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2493 = 7'h25 == _target_predictor_T[6:0] ? 2'h2 : predictor_37; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2494 = 7'h26 == _target_predictor_T[6:0] ? 2'h2 : predictor_38; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2495 = 7'h27 == _target_predictor_T[6:0] ? 2'h2 : predictor_39; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2496 = 7'h28 == _target_predictor_T[6:0] ? 2'h2 : predictor_40; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2497 = 7'h29 == _target_predictor_T[6:0] ? 2'h2 : predictor_41; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2498 = 7'h2a == _target_predictor_T[6:0] ? 2'h2 : predictor_42; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2499 = 7'h2b == _target_predictor_T[6:0] ? 2'h2 : predictor_43; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2500 = 7'h2c == _target_predictor_T[6:0] ? 2'h2 : predictor_44; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2501 = 7'h2d == _target_predictor_T[6:0] ? 2'h2 : predictor_45; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2502 = 7'h2e == _target_predictor_T[6:0] ? 2'h2 : predictor_46; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2503 = 7'h2f == _target_predictor_T[6:0] ? 2'h2 : predictor_47; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2504 = 7'h30 == _target_predictor_T[6:0] ? 2'h2 : predictor_48; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2505 = 7'h31 == _target_predictor_T[6:0] ? 2'h2 : predictor_49; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2506 = 7'h32 == _target_predictor_T[6:0] ? 2'h2 : predictor_50; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2507 = 7'h33 == _target_predictor_T[6:0] ? 2'h2 : predictor_51; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2508 = 7'h34 == _target_predictor_T[6:0] ? 2'h2 : predictor_52; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2509 = 7'h35 == _target_predictor_T[6:0] ? 2'h2 : predictor_53; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2510 = 7'h36 == _target_predictor_T[6:0] ? 2'h2 : predictor_54; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2511 = 7'h37 == _target_predictor_T[6:0] ? 2'h2 : predictor_55; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2512 = 7'h38 == _target_predictor_T[6:0] ? 2'h2 : predictor_56; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2513 = 7'h39 == _target_predictor_T[6:0] ? 2'h2 : predictor_57; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2514 = 7'h3a == _target_predictor_T[6:0] ? 2'h2 : predictor_58; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2515 = 7'h3b == _target_predictor_T[6:0] ? 2'h2 : predictor_59; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2516 = 7'h3c == _target_predictor_T[6:0] ? 2'h2 : predictor_60; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2517 = 7'h3d == _target_predictor_T[6:0] ? 2'h2 : predictor_61; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2518 = 7'h3e == _target_predictor_T[6:0] ? 2'h2 : predictor_62; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2519 = 7'h3f == _target_predictor_T[6:0] ? 2'h2 : predictor_63; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2520 = 7'h40 == _target_predictor_T[6:0] ? 2'h2 : predictor_64; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2521 = 7'h41 == _target_predictor_T[6:0] ? 2'h2 : predictor_65; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2522 = 7'h42 == _target_predictor_T[6:0] ? 2'h2 : predictor_66; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2523 = 7'h43 == _target_predictor_T[6:0] ? 2'h2 : predictor_67; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2524 = 7'h44 == _target_predictor_T[6:0] ? 2'h2 : predictor_68; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2525 = 7'h45 == _target_predictor_T[6:0] ? 2'h2 : predictor_69; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2526 = 7'h46 == _target_predictor_T[6:0] ? 2'h2 : predictor_70; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2527 = 7'h47 == _target_predictor_T[6:0] ? 2'h2 : predictor_71; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2528 = 7'h48 == _target_predictor_T[6:0] ? 2'h2 : predictor_72; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2529 = 7'h49 == _target_predictor_T[6:0] ? 2'h2 : predictor_73; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2530 = 7'h4a == _target_predictor_T[6:0] ? 2'h2 : predictor_74; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2531 = 7'h4b == _target_predictor_T[6:0] ? 2'h2 : predictor_75; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2532 = 7'h4c == _target_predictor_T[6:0] ? 2'h2 : predictor_76; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2533 = 7'h4d == _target_predictor_T[6:0] ? 2'h2 : predictor_77; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2534 = 7'h4e == _target_predictor_T[6:0] ? 2'h2 : predictor_78; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2535 = 7'h4f == _target_predictor_T[6:0] ? 2'h2 : predictor_79; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2536 = 7'h50 == _target_predictor_T[6:0] ? 2'h2 : predictor_80; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2537 = 7'h51 == _target_predictor_T[6:0] ? 2'h2 : predictor_81; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2538 = 7'h52 == _target_predictor_T[6:0] ? 2'h2 : predictor_82; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2539 = 7'h53 == _target_predictor_T[6:0] ? 2'h2 : predictor_83; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2540 = 7'h54 == _target_predictor_T[6:0] ? 2'h2 : predictor_84; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2541 = 7'h55 == _target_predictor_T[6:0] ? 2'h2 : predictor_85; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2542 = 7'h56 == _target_predictor_T[6:0] ? 2'h2 : predictor_86; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2543 = 7'h57 == _target_predictor_T[6:0] ? 2'h2 : predictor_87; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2544 = 7'h58 == _target_predictor_T[6:0] ? 2'h2 : predictor_88; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2545 = 7'h59 == _target_predictor_T[6:0] ? 2'h2 : predictor_89; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2546 = 7'h5a == _target_predictor_T[6:0] ? 2'h2 : predictor_90; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2547 = 7'h5b == _target_predictor_T[6:0] ? 2'h2 : predictor_91; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2548 = 7'h5c == _target_predictor_T[6:0] ? 2'h2 : predictor_92; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2549 = 7'h5d == _target_predictor_T[6:0] ? 2'h2 : predictor_93; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2550 = 7'h5e == _target_predictor_T[6:0] ? 2'h2 : predictor_94; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2551 = 7'h5f == _target_predictor_T[6:0] ? 2'h2 : predictor_95; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2552 = 7'h60 == _target_predictor_T[6:0] ? 2'h2 : predictor_96; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2553 = 7'h61 == _target_predictor_T[6:0] ? 2'h2 : predictor_97; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2554 = 7'h62 == _target_predictor_T[6:0] ? 2'h2 : predictor_98; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2555 = 7'h63 == _target_predictor_T[6:0] ? 2'h2 : predictor_99; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2556 = 7'h64 == _target_predictor_T[6:0] ? 2'h2 : predictor_100; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2557 = 7'h65 == _target_predictor_T[6:0] ? 2'h2 : predictor_101; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2558 = 7'h66 == _target_predictor_T[6:0] ? 2'h2 : predictor_102; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2559 = 7'h67 == _target_predictor_T[6:0] ? 2'h2 : predictor_103; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2560 = 7'h68 == _target_predictor_T[6:0] ? 2'h2 : predictor_104; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2561 = 7'h69 == _target_predictor_T[6:0] ? 2'h2 : predictor_105; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2562 = 7'h6a == _target_predictor_T[6:0] ? 2'h2 : predictor_106; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2563 = 7'h6b == _target_predictor_T[6:0] ? 2'h2 : predictor_107; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2564 = 7'h6c == _target_predictor_T[6:0] ? 2'h2 : predictor_108; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2565 = 7'h6d == _target_predictor_T[6:0] ? 2'h2 : predictor_109; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2566 = 7'h6e == _target_predictor_T[6:0] ? 2'h2 : predictor_110; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2567 = 7'h6f == _target_predictor_T[6:0] ? 2'h2 : predictor_111; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2568 = 7'h70 == _target_predictor_T[6:0] ? 2'h2 : predictor_112; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2569 = 7'h71 == _target_predictor_T[6:0] ? 2'h2 : predictor_113; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2570 = 7'h72 == _target_predictor_T[6:0] ? 2'h2 : predictor_114; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2571 = 7'h73 == _target_predictor_T[6:0] ? 2'h2 : predictor_115; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2572 = 7'h74 == _target_predictor_T[6:0] ? 2'h2 : predictor_116; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2573 = 7'h75 == _target_predictor_T[6:0] ? 2'h2 : predictor_117; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2574 = 7'h76 == _target_predictor_T[6:0] ? 2'h2 : predictor_118; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2575 = 7'h77 == _target_predictor_T[6:0] ? 2'h2 : predictor_119; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2576 = 7'h78 == _target_predictor_T[6:0] ? 2'h2 : predictor_120; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2577 = 7'h79 == _target_predictor_T[6:0] ? 2'h2 : predictor_121; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2578 = 7'h7a == _target_predictor_T[6:0] ? 2'h2 : predictor_122; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2579 = 7'h7b == _target_predictor_T[6:0] ? 2'h2 : predictor_123; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2580 = 7'h7c == _target_predictor_T[6:0] ? 2'h2 : predictor_124; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2581 = 7'h7d == _target_predictor_T[6:0] ? 2'h2 : predictor_125; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2582 = 7'h7e == _target_predictor_T[6:0] ? 2'h2 : predictor_126; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2583 = 7'h7f == _target_predictor_T[6:0] ? 2'h2 : predictor_127; // @[Bpu.scala 154:28 Bpu.scala 154:28 Bpu.scala 74:31]
  wire [1:0] _GEN_2584 = io_branch_info_i_bits_is_taken ? _GEN_1560 : _GEN_2456; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2585 = io_branch_info_i_bits_is_taken ? _GEN_1561 : _GEN_2457; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2586 = io_branch_info_i_bits_is_taken ? _GEN_1562 : _GEN_2458; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2587 = io_branch_info_i_bits_is_taken ? _GEN_1563 : _GEN_2459; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2588 = io_branch_info_i_bits_is_taken ? _GEN_1564 : _GEN_2460; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2589 = io_branch_info_i_bits_is_taken ? _GEN_1565 : _GEN_2461; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2590 = io_branch_info_i_bits_is_taken ? _GEN_1566 : _GEN_2462; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2591 = io_branch_info_i_bits_is_taken ? _GEN_1567 : _GEN_2463; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2592 = io_branch_info_i_bits_is_taken ? _GEN_1568 : _GEN_2464; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2593 = io_branch_info_i_bits_is_taken ? _GEN_1569 : _GEN_2465; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2594 = io_branch_info_i_bits_is_taken ? _GEN_1570 : _GEN_2466; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2595 = io_branch_info_i_bits_is_taken ? _GEN_1571 : _GEN_2467; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2596 = io_branch_info_i_bits_is_taken ? _GEN_1572 : _GEN_2468; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2597 = io_branch_info_i_bits_is_taken ? _GEN_1573 : _GEN_2469; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2598 = io_branch_info_i_bits_is_taken ? _GEN_1574 : _GEN_2470; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2599 = io_branch_info_i_bits_is_taken ? _GEN_1575 : _GEN_2471; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2600 = io_branch_info_i_bits_is_taken ? _GEN_1576 : _GEN_2472; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2601 = io_branch_info_i_bits_is_taken ? _GEN_1577 : _GEN_2473; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2602 = io_branch_info_i_bits_is_taken ? _GEN_1578 : _GEN_2474; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2603 = io_branch_info_i_bits_is_taken ? _GEN_1579 : _GEN_2475; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2604 = io_branch_info_i_bits_is_taken ? _GEN_1580 : _GEN_2476; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2605 = io_branch_info_i_bits_is_taken ? _GEN_1581 : _GEN_2477; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2606 = io_branch_info_i_bits_is_taken ? _GEN_1582 : _GEN_2478; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2607 = io_branch_info_i_bits_is_taken ? _GEN_1583 : _GEN_2479; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2608 = io_branch_info_i_bits_is_taken ? _GEN_1584 : _GEN_2480; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2609 = io_branch_info_i_bits_is_taken ? _GEN_1585 : _GEN_2481; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2610 = io_branch_info_i_bits_is_taken ? _GEN_1586 : _GEN_2482; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2611 = io_branch_info_i_bits_is_taken ? _GEN_1587 : _GEN_2483; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2612 = io_branch_info_i_bits_is_taken ? _GEN_1588 : _GEN_2484; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2613 = io_branch_info_i_bits_is_taken ? _GEN_1589 : _GEN_2485; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2614 = io_branch_info_i_bits_is_taken ? _GEN_1590 : _GEN_2486; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2615 = io_branch_info_i_bits_is_taken ? _GEN_1591 : _GEN_2487; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2616 = io_branch_info_i_bits_is_taken ? _GEN_1592 : _GEN_2488; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2617 = io_branch_info_i_bits_is_taken ? _GEN_1593 : _GEN_2489; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2618 = io_branch_info_i_bits_is_taken ? _GEN_1594 : _GEN_2490; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2619 = io_branch_info_i_bits_is_taken ? _GEN_1595 : _GEN_2491; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2620 = io_branch_info_i_bits_is_taken ? _GEN_1596 : _GEN_2492; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2621 = io_branch_info_i_bits_is_taken ? _GEN_1597 : _GEN_2493; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2622 = io_branch_info_i_bits_is_taken ? _GEN_1598 : _GEN_2494; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2623 = io_branch_info_i_bits_is_taken ? _GEN_1599 : _GEN_2495; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2624 = io_branch_info_i_bits_is_taken ? _GEN_1600 : _GEN_2496; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2625 = io_branch_info_i_bits_is_taken ? _GEN_1601 : _GEN_2497; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2626 = io_branch_info_i_bits_is_taken ? _GEN_1602 : _GEN_2498; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2627 = io_branch_info_i_bits_is_taken ? _GEN_1603 : _GEN_2499; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2628 = io_branch_info_i_bits_is_taken ? _GEN_1604 : _GEN_2500; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2629 = io_branch_info_i_bits_is_taken ? _GEN_1605 : _GEN_2501; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2630 = io_branch_info_i_bits_is_taken ? _GEN_1606 : _GEN_2502; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2631 = io_branch_info_i_bits_is_taken ? _GEN_1607 : _GEN_2503; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2632 = io_branch_info_i_bits_is_taken ? _GEN_1608 : _GEN_2504; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2633 = io_branch_info_i_bits_is_taken ? _GEN_1609 : _GEN_2505; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2634 = io_branch_info_i_bits_is_taken ? _GEN_1610 : _GEN_2506; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2635 = io_branch_info_i_bits_is_taken ? _GEN_1611 : _GEN_2507; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2636 = io_branch_info_i_bits_is_taken ? _GEN_1612 : _GEN_2508; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2637 = io_branch_info_i_bits_is_taken ? _GEN_1613 : _GEN_2509; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2638 = io_branch_info_i_bits_is_taken ? _GEN_1614 : _GEN_2510; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2639 = io_branch_info_i_bits_is_taken ? _GEN_1615 : _GEN_2511; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2640 = io_branch_info_i_bits_is_taken ? _GEN_1616 : _GEN_2512; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2641 = io_branch_info_i_bits_is_taken ? _GEN_1617 : _GEN_2513; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2642 = io_branch_info_i_bits_is_taken ? _GEN_1618 : _GEN_2514; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2643 = io_branch_info_i_bits_is_taken ? _GEN_1619 : _GEN_2515; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2644 = io_branch_info_i_bits_is_taken ? _GEN_1620 : _GEN_2516; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2645 = io_branch_info_i_bits_is_taken ? _GEN_1621 : _GEN_2517; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2646 = io_branch_info_i_bits_is_taken ? _GEN_1622 : _GEN_2518; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2647 = io_branch_info_i_bits_is_taken ? _GEN_1623 : _GEN_2519; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2648 = io_branch_info_i_bits_is_taken ? _GEN_1624 : _GEN_2520; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2649 = io_branch_info_i_bits_is_taken ? _GEN_1625 : _GEN_2521; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2650 = io_branch_info_i_bits_is_taken ? _GEN_1626 : _GEN_2522; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2651 = io_branch_info_i_bits_is_taken ? _GEN_1627 : _GEN_2523; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2652 = io_branch_info_i_bits_is_taken ? _GEN_1628 : _GEN_2524; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2653 = io_branch_info_i_bits_is_taken ? _GEN_1629 : _GEN_2525; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2654 = io_branch_info_i_bits_is_taken ? _GEN_1630 : _GEN_2526; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2655 = io_branch_info_i_bits_is_taken ? _GEN_1631 : _GEN_2527; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2656 = io_branch_info_i_bits_is_taken ? _GEN_1632 : _GEN_2528; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2657 = io_branch_info_i_bits_is_taken ? _GEN_1633 : _GEN_2529; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2658 = io_branch_info_i_bits_is_taken ? _GEN_1634 : _GEN_2530; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2659 = io_branch_info_i_bits_is_taken ? _GEN_1635 : _GEN_2531; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2660 = io_branch_info_i_bits_is_taken ? _GEN_1636 : _GEN_2532; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2661 = io_branch_info_i_bits_is_taken ? _GEN_1637 : _GEN_2533; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2662 = io_branch_info_i_bits_is_taken ? _GEN_1638 : _GEN_2534; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2663 = io_branch_info_i_bits_is_taken ? _GEN_1639 : _GEN_2535; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2664 = io_branch_info_i_bits_is_taken ? _GEN_1640 : _GEN_2536; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2665 = io_branch_info_i_bits_is_taken ? _GEN_1641 : _GEN_2537; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2666 = io_branch_info_i_bits_is_taken ? _GEN_1642 : _GEN_2538; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2667 = io_branch_info_i_bits_is_taken ? _GEN_1643 : _GEN_2539; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2668 = io_branch_info_i_bits_is_taken ? _GEN_1644 : _GEN_2540; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2669 = io_branch_info_i_bits_is_taken ? _GEN_1645 : _GEN_2541; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2670 = io_branch_info_i_bits_is_taken ? _GEN_1646 : _GEN_2542; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2671 = io_branch_info_i_bits_is_taken ? _GEN_1647 : _GEN_2543; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2672 = io_branch_info_i_bits_is_taken ? _GEN_1648 : _GEN_2544; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2673 = io_branch_info_i_bits_is_taken ? _GEN_1649 : _GEN_2545; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2674 = io_branch_info_i_bits_is_taken ? _GEN_1650 : _GEN_2546; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2675 = io_branch_info_i_bits_is_taken ? _GEN_1651 : _GEN_2547; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2676 = io_branch_info_i_bits_is_taken ? _GEN_1652 : _GEN_2548; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2677 = io_branch_info_i_bits_is_taken ? _GEN_1653 : _GEN_2549; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2678 = io_branch_info_i_bits_is_taken ? _GEN_1654 : _GEN_2550; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2679 = io_branch_info_i_bits_is_taken ? _GEN_1655 : _GEN_2551; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2680 = io_branch_info_i_bits_is_taken ? _GEN_1656 : _GEN_2552; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2681 = io_branch_info_i_bits_is_taken ? _GEN_1657 : _GEN_2553; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2682 = io_branch_info_i_bits_is_taken ? _GEN_1658 : _GEN_2554; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2683 = io_branch_info_i_bits_is_taken ? _GEN_1659 : _GEN_2555; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2684 = io_branch_info_i_bits_is_taken ? _GEN_1660 : _GEN_2556; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2685 = io_branch_info_i_bits_is_taken ? _GEN_1661 : _GEN_2557; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2686 = io_branch_info_i_bits_is_taken ? _GEN_1662 : _GEN_2558; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2687 = io_branch_info_i_bits_is_taken ? _GEN_1663 : _GEN_2559; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2688 = io_branch_info_i_bits_is_taken ? _GEN_1664 : _GEN_2560; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2689 = io_branch_info_i_bits_is_taken ? _GEN_1665 : _GEN_2561; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2690 = io_branch_info_i_bits_is_taken ? _GEN_1666 : _GEN_2562; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2691 = io_branch_info_i_bits_is_taken ? _GEN_1667 : _GEN_2563; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2692 = io_branch_info_i_bits_is_taken ? _GEN_1668 : _GEN_2564; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2693 = io_branch_info_i_bits_is_taken ? _GEN_1669 : _GEN_2565; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2694 = io_branch_info_i_bits_is_taken ? _GEN_1670 : _GEN_2566; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2695 = io_branch_info_i_bits_is_taken ? _GEN_1671 : _GEN_2567; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2696 = io_branch_info_i_bits_is_taken ? _GEN_1672 : _GEN_2568; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2697 = io_branch_info_i_bits_is_taken ? _GEN_1673 : _GEN_2569; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2698 = io_branch_info_i_bits_is_taken ? _GEN_1674 : _GEN_2570; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2699 = io_branch_info_i_bits_is_taken ? _GEN_1675 : _GEN_2571; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2700 = io_branch_info_i_bits_is_taken ? _GEN_1676 : _GEN_2572; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2701 = io_branch_info_i_bits_is_taken ? _GEN_1677 : _GEN_2573; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2702 = io_branch_info_i_bits_is_taken ? _GEN_1678 : _GEN_2574; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2703 = io_branch_info_i_bits_is_taken ? _GEN_1679 : _GEN_2575; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2704 = io_branch_info_i_bits_is_taken ? _GEN_1680 : _GEN_2576; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2705 = io_branch_info_i_bits_is_taken ? _GEN_1681 : _GEN_2577; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2706 = io_branch_info_i_bits_is_taken ? _GEN_1682 : _GEN_2578; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2707 = io_branch_info_i_bits_is_taken ? _GEN_1683 : _GEN_2579; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2708 = io_branch_info_i_bits_is_taken ? _GEN_1684 : _GEN_2580; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2709 = io_branch_info_i_bits_is_taken ? _GEN_1685 : _GEN_2581; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2710 = io_branch_info_i_bits_is_taken ? _GEN_1686 : _GEN_2582; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2711 = io_branch_info_i_bits_is_taken ? _GEN_1687 : _GEN_2583; // @[Bpu.scala 151:46]
  wire [1:0] _GEN_2712 = _T_6 ? _GEN_2584 : predictor_0; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2713 = _T_6 ? _GEN_2585 : predictor_1; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2714 = _T_6 ? _GEN_2586 : predictor_2; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2715 = _T_6 ? _GEN_2587 : predictor_3; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2716 = _T_6 ? _GEN_2588 : predictor_4; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2717 = _T_6 ? _GEN_2589 : predictor_5; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2718 = _T_6 ? _GEN_2590 : predictor_6; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2719 = _T_6 ? _GEN_2591 : predictor_7; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2720 = _T_6 ? _GEN_2592 : predictor_8; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2721 = _T_6 ? _GEN_2593 : predictor_9; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2722 = _T_6 ? _GEN_2594 : predictor_10; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2723 = _T_6 ? _GEN_2595 : predictor_11; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2724 = _T_6 ? _GEN_2596 : predictor_12; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2725 = _T_6 ? _GEN_2597 : predictor_13; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2726 = _T_6 ? _GEN_2598 : predictor_14; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2727 = _T_6 ? _GEN_2599 : predictor_15; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2728 = _T_6 ? _GEN_2600 : predictor_16; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2729 = _T_6 ? _GEN_2601 : predictor_17; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2730 = _T_6 ? _GEN_2602 : predictor_18; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2731 = _T_6 ? _GEN_2603 : predictor_19; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2732 = _T_6 ? _GEN_2604 : predictor_20; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2733 = _T_6 ? _GEN_2605 : predictor_21; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2734 = _T_6 ? _GEN_2606 : predictor_22; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2735 = _T_6 ? _GEN_2607 : predictor_23; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2736 = _T_6 ? _GEN_2608 : predictor_24; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2737 = _T_6 ? _GEN_2609 : predictor_25; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2738 = _T_6 ? _GEN_2610 : predictor_26; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2739 = _T_6 ? _GEN_2611 : predictor_27; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2740 = _T_6 ? _GEN_2612 : predictor_28; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2741 = _T_6 ? _GEN_2613 : predictor_29; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2742 = _T_6 ? _GEN_2614 : predictor_30; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2743 = _T_6 ? _GEN_2615 : predictor_31; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2744 = _T_6 ? _GEN_2616 : predictor_32; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2745 = _T_6 ? _GEN_2617 : predictor_33; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2746 = _T_6 ? _GEN_2618 : predictor_34; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2747 = _T_6 ? _GEN_2619 : predictor_35; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2748 = _T_6 ? _GEN_2620 : predictor_36; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2749 = _T_6 ? _GEN_2621 : predictor_37; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2750 = _T_6 ? _GEN_2622 : predictor_38; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2751 = _T_6 ? _GEN_2623 : predictor_39; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2752 = _T_6 ? _GEN_2624 : predictor_40; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2753 = _T_6 ? _GEN_2625 : predictor_41; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2754 = _T_6 ? _GEN_2626 : predictor_42; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2755 = _T_6 ? _GEN_2627 : predictor_43; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2756 = _T_6 ? _GEN_2628 : predictor_44; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2757 = _T_6 ? _GEN_2629 : predictor_45; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2758 = _T_6 ? _GEN_2630 : predictor_46; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2759 = _T_6 ? _GEN_2631 : predictor_47; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2760 = _T_6 ? _GEN_2632 : predictor_48; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2761 = _T_6 ? _GEN_2633 : predictor_49; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2762 = _T_6 ? _GEN_2634 : predictor_50; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2763 = _T_6 ? _GEN_2635 : predictor_51; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2764 = _T_6 ? _GEN_2636 : predictor_52; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2765 = _T_6 ? _GEN_2637 : predictor_53; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2766 = _T_6 ? _GEN_2638 : predictor_54; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2767 = _T_6 ? _GEN_2639 : predictor_55; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2768 = _T_6 ? _GEN_2640 : predictor_56; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2769 = _T_6 ? _GEN_2641 : predictor_57; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2770 = _T_6 ? _GEN_2642 : predictor_58; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2771 = _T_6 ? _GEN_2643 : predictor_59; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2772 = _T_6 ? _GEN_2644 : predictor_60; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2773 = _T_6 ? _GEN_2645 : predictor_61; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2774 = _T_6 ? _GEN_2646 : predictor_62; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2775 = _T_6 ? _GEN_2647 : predictor_63; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2776 = _T_6 ? _GEN_2648 : predictor_64; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2777 = _T_6 ? _GEN_2649 : predictor_65; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2778 = _T_6 ? _GEN_2650 : predictor_66; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2779 = _T_6 ? _GEN_2651 : predictor_67; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2780 = _T_6 ? _GEN_2652 : predictor_68; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2781 = _T_6 ? _GEN_2653 : predictor_69; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2782 = _T_6 ? _GEN_2654 : predictor_70; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2783 = _T_6 ? _GEN_2655 : predictor_71; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2784 = _T_6 ? _GEN_2656 : predictor_72; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2785 = _T_6 ? _GEN_2657 : predictor_73; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2786 = _T_6 ? _GEN_2658 : predictor_74; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2787 = _T_6 ? _GEN_2659 : predictor_75; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2788 = _T_6 ? _GEN_2660 : predictor_76; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2789 = _T_6 ? _GEN_2661 : predictor_77; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2790 = _T_6 ? _GEN_2662 : predictor_78; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2791 = _T_6 ? _GEN_2663 : predictor_79; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2792 = _T_6 ? _GEN_2664 : predictor_80; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2793 = _T_6 ? _GEN_2665 : predictor_81; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2794 = _T_6 ? _GEN_2666 : predictor_82; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2795 = _T_6 ? _GEN_2667 : predictor_83; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2796 = _T_6 ? _GEN_2668 : predictor_84; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2797 = _T_6 ? _GEN_2669 : predictor_85; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2798 = _T_6 ? _GEN_2670 : predictor_86; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2799 = _T_6 ? _GEN_2671 : predictor_87; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2800 = _T_6 ? _GEN_2672 : predictor_88; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2801 = _T_6 ? _GEN_2673 : predictor_89; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2802 = _T_6 ? _GEN_2674 : predictor_90; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2803 = _T_6 ? _GEN_2675 : predictor_91; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2804 = _T_6 ? _GEN_2676 : predictor_92; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2805 = _T_6 ? _GEN_2677 : predictor_93; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2806 = _T_6 ? _GEN_2678 : predictor_94; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2807 = _T_6 ? _GEN_2679 : predictor_95; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2808 = _T_6 ? _GEN_2680 : predictor_96; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2809 = _T_6 ? _GEN_2681 : predictor_97; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2810 = _T_6 ? _GEN_2682 : predictor_98; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2811 = _T_6 ? _GEN_2683 : predictor_99; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2812 = _T_6 ? _GEN_2684 : predictor_100; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2813 = _T_6 ? _GEN_2685 : predictor_101; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2814 = _T_6 ? _GEN_2686 : predictor_102; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2815 = _T_6 ? _GEN_2687 : predictor_103; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2816 = _T_6 ? _GEN_2688 : predictor_104; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2817 = _T_6 ? _GEN_2689 : predictor_105; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2818 = _T_6 ? _GEN_2690 : predictor_106; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2819 = _T_6 ? _GEN_2691 : predictor_107; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2820 = _T_6 ? _GEN_2692 : predictor_108; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2821 = _T_6 ? _GEN_2693 : predictor_109; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2822 = _T_6 ? _GEN_2694 : predictor_110; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2823 = _T_6 ? _GEN_2695 : predictor_111; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2824 = _T_6 ? _GEN_2696 : predictor_112; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2825 = _T_6 ? _GEN_2697 : predictor_113; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2826 = _T_6 ? _GEN_2698 : predictor_114; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2827 = _T_6 ? _GEN_2699 : predictor_115; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2828 = _T_6 ? _GEN_2700 : predictor_116; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2829 = _T_6 ? _GEN_2701 : predictor_117; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2830 = _T_6 ? _GEN_2702 : predictor_118; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2831 = _T_6 ? _GEN_2703 : predictor_119; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2832 = _T_6 ? _GEN_2704 : predictor_120; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2833 = _T_6 ? _GEN_2705 : predictor_121; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2834 = _T_6 ? _GEN_2706 : predictor_122; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2835 = _T_6 ? _GEN_2707 : predictor_123; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2836 = _T_6 ? _GEN_2708 : predictor_124; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2837 = _T_6 ? _GEN_2709 : predictor_125; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2838 = _T_6 ? _GEN_2710 : predictor_126; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2839 = _T_6 ? _GEN_2711 : predictor_127; // @[Conditional.scala 39:67 Bpu.scala 74:31]
  wire [1:0] _GEN_2840 = _T_5 ? _GEN_1816 : _GEN_2712; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2841 = _T_5 ? _GEN_1817 : _GEN_2713; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2842 = _T_5 ? _GEN_1818 : _GEN_2714; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2843 = _T_5 ? _GEN_1819 : _GEN_2715; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2844 = _T_5 ? _GEN_1820 : _GEN_2716; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2845 = _T_5 ? _GEN_1821 : _GEN_2717; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2846 = _T_5 ? _GEN_1822 : _GEN_2718; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2847 = _T_5 ? _GEN_1823 : _GEN_2719; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2848 = _T_5 ? _GEN_1824 : _GEN_2720; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2849 = _T_5 ? _GEN_1825 : _GEN_2721; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2850 = _T_5 ? _GEN_1826 : _GEN_2722; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2851 = _T_5 ? _GEN_1827 : _GEN_2723; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2852 = _T_5 ? _GEN_1828 : _GEN_2724; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2853 = _T_5 ? _GEN_1829 : _GEN_2725; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2854 = _T_5 ? _GEN_1830 : _GEN_2726; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2855 = _T_5 ? _GEN_1831 : _GEN_2727; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2856 = _T_5 ? _GEN_1832 : _GEN_2728; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2857 = _T_5 ? _GEN_1833 : _GEN_2729; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2858 = _T_5 ? _GEN_1834 : _GEN_2730; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2859 = _T_5 ? _GEN_1835 : _GEN_2731; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2860 = _T_5 ? _GEN_1836 : _GEN_2732; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2861 = _T_5 ? _GEN_1837 : _GEN_2733; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2862 = _T_5 ? _GEN_1838 : _GEN_2734; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2863 = _T_5 ? _GEN_1839 : _GEN_2735; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2864 = _T_5 ? _GEN_1840 : _GEN_2736; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2865 = _T_5 ? _GEN_1841 : _GEN_2737; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2866 = _T_5 ? _GEN_1842 : _GEN_2738; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2867 = _T_5 ? _GEN_1843 : _GEN_2739; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2868 = _T_5 ? _GEN_1844 : _GEN_2740; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2869 = _T_5 ? _GEN_1845 : _GEN_2741; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2870 = _T_5 ? _GEN_1846 : _GEN_2742; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2871 = _T_5 ? _GEN_1847 : _GEN_2743; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2872 = _T_5 ? _GEN_1848 : _GEN_2744; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2873 = _T_5 ? _GEN_1849 : _GEN_2745; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2874 = _T_5 ? _GEN_1850 : _GEN_2746; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2875 = _T_5 ? _GEN_1851 : _GEN_2747; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2876 = _T_5 ? _GEN_1852 : _GEN_2748; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2877 = _T_5 ? _GEN_1853 : _GEN_2749; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2878 = _T_5 ? _GEN_1854 : _GEN_2750; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2879 = _T_5 ? _GEN_1855 : _GEN_2751; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2880 = _T_5 ? _GEN_1856 : _GEN_2752; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2881 = _T_5 ? _GEN_1857 : _GEN_2753; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2882 = _T_5 ? _GEN_1858 : _GEN_2754; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2883 = _T_5 ? _GEN_1859 : _GEN_2755; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2884 = _T_5 ? _GEN_1860 : _GEN_2756; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2885 = _T_5 ? _GEN_1861 : _GEN_2757; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2886 = _T_5 ? _GEN_1862 : _GEN_2758; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2887 = _T_5 ? _GEN_1863 : _GEN_2759; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2888 = _T_5 ? _GEN_1864 : _GEN_2760; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2889 = _T_5 ? _GEN_1865 : _GEN_2761; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2890 = _T_5 ? _GEN_1866 : _GEN_2762; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2891 = _T_5 ? _GEN_1867 : _GEN_2763; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2892 = _T_5 ? _GEN_1868 : _GEN_2764; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2893 = _T_5 ? _GEN_1869 : _GEN_2765; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2894 = _T_5 ? _GEN_1870 : _GEN_2766; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2895 = _T_5 ? _GEN_1871 : _GEN_2767; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2896 = _T_5 ? _GEN_1872 : _GEN_2768; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2897 = _T_5 ? _GEN_1873 : _GEN_2769; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2898 = _T_5 ? _GEN_1874 : _GEN_2770; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2899 = _T_5 ? _GEN_1875 : _GEN_2771; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2900 = _T_5 ? _GEN_1876 : _GEN_2772; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2901 = _T_5 ? _GEN_1877 : _GEN_2773; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2902 = _T_5 ? _GEN_1878 : _GEN_2774; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2903 = _T_5 ? _GEN_1879 : _GEN_2775; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2904 = _T_5 ? _GEN_1880 : _GEN_2776; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2905 = _T_5 ? _GEN_1881 : _GEN_2777; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2906 = _T_5 ? _GEN_1882 : _GEN_2778; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2907 = _T_5 ? _GEN_1883 : _GEN_2779; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2908 = _T_5 ? _GEN_1884 : _GEN_2780; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2909 = _T_5 ? _GEN_1885 : _GEN_2781; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2910 = _T_5 ? _GEN_1886 : _GEN_2782; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2911 = _T_5 ? _GEN_1887 : _GEN_2783; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2912 = _T_5 ? _GEN_1888 : _GEN_2784; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2913 = _T_5 ? _GEN_1889 : _GEN_2785; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2914 = _T_5 ? _GEN_1890 : _GEN_2786; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2915 = _T_5 ? _GEN_1891 : _GEN_2787; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2916 = _T_5 ? _GEN_1892 : _GEN_2788; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2917 = _T_5 ? _GEN_1893 : _GEN_2789; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2918 = _T_5 ? _GEN_1894 : _GEN_2790; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2919 = _T_5 ? _GEN_1895 : _GEN_2791; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2920 = _T_5 ? _GEN_1896 : _GEN_2792; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2921 = _T_5 ? _GEN_1897 : _GEN_2793; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2922 = _T_5 ? _GEN_1898 : _GEN_2794; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2923 = _T_5 ? _GEN_1899 : _GEN_2795; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2924 = _T_5 ? _GEN_1900 : _GEN_2796; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2925 = _T_5 ? _GEN_1901 : _GEN_2797; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2926 = _T_5 ? _GEN_1902 : _GEN_2798; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2927 = _T_5 ? _GEN_1903 : _GEN_2799; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2928 = _T_5 ? _GEN_1904 : _GEN_2800; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2929 = _T_5 ? _GEN_1905 : _GEN_2801; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2930 = _T_5 ? _GEN_1906 : _GEN_2802; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2931 = _T_5 ? _GEN_1907 : _GEN_2803; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2932 = _T_5 ? _GEN_1908 : _GEN_2804; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2933 = _T_5 ? _GEN_1909 : _GEN_2805; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2934 = _T_5 ? _GEN_1910 : _GEN_2806; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2935 = _T_5 ? _GEN_1911 : _GEN_2807; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2936 = _T_5 ? _GEN_1912 : _GEN_2808; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2937 = _T_5 ? _GEN_1913 : _GEN_2809; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2938 = _T_5 ? _GEN_1914 : _GEN_2810; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2939 = _T_5 ? _GEN_1915 : _GEN_2811; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2940 = _T_5 ? _GEN_1916 : _GEN_2812; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2941 = _T_5 ? _GEN_1917 : _GEN_2813; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2942 = _T_5 ? _GEN_1918 : _GEN_2814; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2943 = _T_5 ? _GEN_1919 : _GEN_2815; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2944 = _T_5 ? _GEN_1920 : _GEN_2816; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2945 = _T_5 ? _GEN_1921 : _GEN_2817; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2946 = _T_5 ? _GEN_1922 : _GEN_2818; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2947 = _T_5 ? _GEN_1923 : _GEN_2819; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2948 = _T_5 ? _GEN_1924 : _GEN_2820; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2949 = _T_5 ? _GEN_1925 : _GEN_2821; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2950 = _T_5 ? _GEN_1926 : _GEN_2822; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2951 = _T_5 ? _GEN_1927 : _GEN_2823; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2952 = _T_5 ? _GEN_1928 : _GEN_2824; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2953 = _T_5 ? _GEN_1929 : _GEN_2825; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2954 = _T_5 ? _GEN_1930 : _GEN_2826; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2955 = _T_5 ? _GEN_1931 : _GEN_2827; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2956 = _T_5 ? _GEN_1932 : _GEN_2828; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2957 = _T_5 ? _GEN_1933 : _GEN_2829; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2958 = _T_5 ? _GEN_1934 : _GEN_2830; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2959 = _T_5 ? _GEN_1935 : _GEN_2831; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2960 = _T_5 ? _GEN_1936 : _GEN_2832; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2961 = _T_5 ? _GEN_1937 : _GEN_2833; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2962 = _T_5 ? _GEN_1938 : _GEN_2834; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2963 = _T_5 ? _GEN_1939 : _GEN_2835; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2964 = _T_5 ? _GEN_1940 : _GEN_2836; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2965 = _T_5 ? _GEN_1941 : _GEN_2837; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2966 = _T_5 ? _GEN_1942 : _GEN_2838; // @[Conditional.scala 39:67]
  wire [1:0] _GEN_2967 = _T_5 ? _GEN_1943 : _GEN_2839; // @[Conditional.scala 39:67]
  reg [31:0] bpu_inst_packet_o_data_0; // @[Bpu.scala 165:30]
  reg [31:0] bpu_inst_packet_o_data_1; // @[Bpu.scala 165:30]
  reg [31:0] bpu_inst_packet_o_data_2; // @[Bpu.scala 165:30]
  reg [31:0] bpu_inst_packet_o_data_3; // @[Bpu.scala 165:30]
  reg [31:0] bpu_inst_packet_o_data_4; // @[Bpu.scala 165:30]
  reg [31:0] bpu_inst_packet_o_data_5; // @[Bpu.scala 165:30]
  reg [31:0] bpu_inst_packet_o_data_6; // @[Bpu.scala 165:30]
  reg [31:0] bpu_inst_packet_o_data_7; // @[Bpu.scala 165:30]
  reg [31:0] bpu_inst_packet_o_addr; // @[Bpu.scala 165:30]
  reg [3:0] bpu_inst_packet_o_gh_backup; // @[Bpu.scala 165:30]
  reg  bpu_inst_packet_o_valid_mask_0; // @[Bpu.scala 165:30]
  reg  bpu_inst_packet_o_valid_mask_1; // @[Bpu.scala 165:30]
  reg  bpu_inst_packet_o_valid_mask_2; // @[Bpu.scala 165:30]
  reg  bpu_inst_packet_o_valid_mask_3; // @[Bpu.scala 165:30]
  reg  bpu_inst_packet_o_valid_mask_4; // @[Bpu.scala 165:30]
  reg  bpu_inst_packet_o_valid_mask_5; // @[Bpu.scala 165:30]
  reg  bpu_inst_packet_o_valid_mask_6; // @[Bpu.scala 165:30]
  reg  bpu_inst_packet_o_valid_mask_7; // @[Bpu.scala 165:30]
  reg  bpu_inst_packet_o_predict_mask_0; // @[Bpu.scala 165:30]
  reg  bpu_inst_packet_o_predict_mask_1; // @[Bpu.scala 165:30]
  reg  bpu_inst_packet_o_predict_mask_2; // @[Bpu.scala 165:30]
  reg  bpu_inst_packet_o_predict_mask_3; // @[Bpu.scala 165:30]
  reg  bpu_inst_packet_o_predict_mask_4; // @[Bpu.scala 165:30]
  reg  bpu_inst_packet_o_predict_mask_5; // @[Bpu.scala 165:30]
  reg  bpu_inst_packet_o_predict_mask_6; // @[Bpu.scala 165:30]
  reg  bpu_inst_packet_o_predict_mask_7; // @[Bpu.scala 165:30]
  reg  bpu_inst_packet_o_valid; // @[Bpu.scala 166:40]
  wire [3:0] io_bpu_debug_branch_mask_lo = {branch_mask_3,branch_mask_2,branch_mask_1,branch_mask_0}; // @[Bpu.scala 201:56]
  wire [3:0] io_bpu_debug_branch_mask_hi = {branch_mask_7,branch_mask_6,branch_mask_5,branch_mask_4}; // @[Bpu.scala 201:56]
  wire [3:0] io_bpu_debug_fetched_mask_lo = {fetched_mask_3,fetched_mask_2,fetched_mask_1,fetched_mask_0}; // @[Bpu.scala 202:58]
  wire [3:0] io_bpu_debug_fetched_mask_hi = {fetched_mask_7,fetched_mask_6,fetched_mask_5,fetched_mask_4}; // @[Bpu.scala 202:58]
  assign io_resp_o_valid = io_inst_packet_i_valid; // @[Bpu.scala 163:19]
  assign io_resp_o_bits_predict_addr = $signed(_predict_addr_T_5) + 32'sh4; // @[Bpu.scala 110:145]
  assign io_resp_o_bits_is_taken = |_is_taken_T; // @[Bpu.scala 100:54]
  assign io_resp_o_bits_take_delay = inst_idx == 3'h7 & is_taken; // @[Bpu.scala 117:53]
  assign io_bpu_inst_packet_o_valid = bpu_inst_packet_o_valid; // @[Bpu.scala 179:29]
  assign io_bpu_inst_packet_o_bits_data_0 = bpu_inst_packet_o_data_0; // @[Bpu.scala 178:28]
  assign io_bpu_inst_packet_o_bits_data_1 = bpu_inst_packet_o_data_1; // @[Bpu.scala 178:28]
  assign io_bpu_inst_packet_o_bits_data_2 = bpu_inst_packet_o_data_2; // @[Bpu.scala 178:28]
  assign io_bpu_inst_packet_o_bits_data_3 = bpu_inst_packet_o_data_3; // @[Bpu.scala 178:28]
  assign io_bpu_inst_packet_o_bits_data_4 = bpu_inst_packet_o_data_4; // @[Bpu.scala 178:28]
  assign io_bpu_inst_packet_o_bits_data_5 = bpu_inst_packet_o_data_5; // @[Bpu.scala 178:28]
  assign io_bpu_inst_packet_o_bits_data_6 = bpu_inst_packet_o_data_6; // @[Bpu.scala 178:28]
  assign io_bpu_inst_packet_o_bits_data_7 = bpu_inst_packet_o_data_7; // @[Bpu.scala 178:28]
  assign io_bpu_inst_packet_o_bits_addr = bpu_inst_packet_o_addr; // @[Bpu.scala 178:28]
  assign io_bpu_inst_packet_o_bits_gh_backup = bpu_inst_packet_o_gh_backup; // @[Bpu.scala 178:28]
  assign io_bpu_inst_packet_o_bits_valid_mask_0 = bpu_inst_packet_o_valid_mask_0; // @[Bpu.scala 178:28]
  assign io_bpu_inst_packet_o_bits_valid_mask_1 = bpu_inst_packet_o_valid_mask_1; // @[Bpu.scala 178:28]
  assign io_bpu_inst_packet_o_bits_valid_mask_2 = bpu_inst_packet_o_valid_mask_2; // @[Bpu.scala 178:28]
  assign io_bpu_inst_packet_o_bits_valid_mask_3 = bpu_inst_packet_o_valid_mask_3; // @[Bpu.scala 178:28]
  assign io_bpu_inst_packet_o_bits_valid_mask_4 = bpu_inst_packet_o_valid_mask_4; // @[Bpu.scala 178:28]
  assign io_bpu_inst_packet_o_bits_valid_mask_5 = bpu_inst_packet_o_valid_mask_5; // @[Bpu.scala 178:28]
  assign io_bpu_inst_packet_o_bits_valid_mask_6 = bpu_inst_packet_o_valid_mask_6; // @[Bpu.scala 178:28]
  assign io_bpu_inst_packet_o_bits_valid_mask_7 = bpu_inst_packet_o_valid_mask_7; // @[Bpu.scala 178:28]
  assign io_bpu_inst_packet_o_bits_predict_mask_0 = bpu_inst_packet_o_predict_mask_0; // @[Bpu.scala 178:28]
  assign io_bpu_inst_packet_o_bits_predict_mask_1 = bpu_inst_packet_o_predict_mask_1; // @[Bpu.scala 178:28]
  assign io_bpu_inst_packet_o_bits_predict_mask_2 = bpu_inst_packet_o_predict_mask_2; // @[Bpu.scala 178:28]
  assign io_bpu_inst_packet_o_bits_predict_mask_3 = bpu_inst_packet_o_predict_mask_3; // @[Bpu.scala 178:28]
  assign io_bpu_inst_packet_o_bits_predict_mask_4 = bpu_inst_packet_o_predict_mask_4; // @[Bpu.scala 178:28]
  assign io_bpu_inst_packet_o_bits_predict_mask_5 = bpu_inst_packet_o_predict_mask_5; // @[Bpu.scala 178:28]
  assign io_bpu_inst_packet_o_bits_predict_mask_6 = bpu_inst_packet_o_predict_mask_6; // @[Bpu.scala 178:28]
  assign io_bpu_inst_packet_o_bits_predict_mask_7 = bpu_inst_packet_o_predict_mask_7; // @[Bpu.scala 178:28]
  assign io_bpu_debug_branch_mask = {io_bpu_debug_branch_mask_hi,io_bpu_debug_branch_mask_lo}; // @[Bpu.scala 201:56]
  assign io_bpu_debug_fetched_mask = {io_bpu_debug_fetched_mask_hi,io_bpu_debug_fetched_mask_lo}; // @[Bpu.scala 202:58]
  assign io_bpu_debug_predict_branch = {is_taken_hi,is_taken_lo}; // @[Bpu.scala 203:62]
  assign io_bpu_debug_predict_addr = $signed(_predict_addr_T_5) + 32'sh4; // @[Bpu.scala 110:145]
  assign io_bpu_debug_is_taken = |_is_taken_T; // @[Bpu.scala 100:54]
  assign io_bpu_debug_take_delay = inst_idx == 3'h7 & is_taken; // @[Bpu.scala 117:53]
  assign io_bpu_debug_inst_packet_0 = io_inst_packet_i_bits_data_0; // @[Bpu.scala 207:27]
  assign io_bpu_debug_inst_packet_1 = io_inst_packet_i_bits_data_1; // @[Bpu.scala 207:27]
  assign io_bpu_debug_inst_packet_2 = io_inst_packet_i_bits_data_2; // @[Bpu.scala 207:27]
  assign io_bpu_debug_inst_packet_3 = io_inst_packet_i_bits_data_3; // @[Bpu.scala 207:27]
  assign io_bpu_debug_inst_packet_4 = io_inst_packet_i_bits_data_4; // @[Bpu.scala 207:27]
  assign io_bpu_debug_inst_packet_5 = io_inst_packet_i_bits_data_5; // @[Bpu.scala 207:27]
  assign io_bpu_debug_inst_packet_6 = io_inst_packet_i_bits_data_6; // @[Bpu.scala 207:27]
  assign io_bpu_debug_inst_packet_7 = io_inst_packet_i_bits_data_7; // @[Bpu.scala 207:27]
  always @(posedge clock) begin
    if (reset) begin // @[Bpu.scala 73:31]
      global_history <= 4'h0; // @[Bpu.scala 73:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_predict_miss) begin // @[Bpu.scala 125:24]
      global_history <= io_branch_info_i_bits_gh_update;
    end else begin
      global_history <= _hi_T_1;
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_0 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_0 <= _GEN_1176;
        end else begin
          predictor_0 <= _GEN_1304;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_0 <= _GEN_1816;
      end else begin
        predictor_0 <= _GEN_2840;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_1 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_1 <= _GEN_1177;
        end else begin
          predictor_1 <= _GEN_1305;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_1 <= _GEN_1817;
      end else begin
        predictor_1 <= _GEN_2841;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_2 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_2 <= _GEN_1178;
        end else begin
          predictor_2 <= _GEN_1306;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_2 <= _GEN_1818;
      end else begin
        predictor_2 <= _GEN_2842;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_3 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_3 <= _GEN_1179;
        end else begin
          predictor_3 <= _GEN_1307;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_3 <= _GEN_1819;
      end else begin
        predictor_3 <= _GEN_2843;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_4 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_4 <= _GEN_1180;
        end else begin
          predictor_4 <= _GEN_1308;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_4 <= _GEN_1820;
      end else begin
        predictor_4 <= _GEN_2844;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_5 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_5 <= _GEN_1181;
        end else begin
          predictor_5 <= _GEN_1309;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_5 <= _GEN_1821;
      end else begin
        predictor_5 <= _GEN_2845;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_6 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_6 <= _GEN_1182;
        end else begin
          predictor_6 <= _GEN_1310;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_6 <= _GEN_1822;
      end else begin
        predictor_6 <= _GEN_2846;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_7 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_7 <= _GEN_1183;
        end else begin
          predictor_7 <= _GEN_1311;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_7 <= _GEN_1823;
      end else begin
        predictor_7 <= _GEN_2847;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_8 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_8 <= _GEN_1184;
        end else begin
          predictor_8 <= _GEN_1312;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_8 <= _GEN_1824;
      end else begin
        predictor_8 <= _GEN_2848;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_9 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_9 <= _GEN_1185;
        end else begin
          predictor_9 <= _GEN_1313;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_9 <= _GEN_1825;
      end else begin
        predictor_9 <= _GEN_2849;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_10 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_10 <= _GEN_1186;
        end else begin
          predictor_10 <= _GEN_1314;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_10 <= _GEN_1826;
      end else begin
        predictor_10 <= _GEN_2850;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_11 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_11 <= _GEN_1187;
        end else begin
          predictor_11 <= _GEN_1315;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_11 <= _GEN_1827;
      end else begin
        predictor_11 <= _GEN_2851;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_12 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_12 <= _GEN_1188;
        end else begin
          predictor_12 <= _GEN_1316;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_12 <= _GEN_1828;
      end else begin
        predictor_12 <= _GEN_2852;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_13 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_13 <= _GEN_1189;
        end else begin
          predictor_13 <= _GEN_1317;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_13 <= _GEN_1829;
      end else begin
        predictor_13 <= _GEN_2853;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_14 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_14 <= _GEN_1190;
        end else begin
          predictor_14 <= _GEN_1318;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_14 <= _GEN_1830;
      end else begin
        predictor_14 <= _GEN_2854;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_15 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_15 <= _GEN_1191;
        end else begin
          predictor_15 <= _GEN_1319;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_15 <= _GEN_1831;
      end else begin
        predictor_15 <= _GEN_2855;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_16 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_16 <= _GEN_1192;
        end else begin
          predictor_16 <= _GEN_1320;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_16 <= _GEN_1832;
      end else begin
        predictor_16 <= _GEN_2856;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_17 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_17 <= _GEN_1193;
        end else begin
          predictor_17 <= _GEN_1321;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_17 <= _GEN_1833;
      end else begin
        predictor_17 <= _GEN_2857;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_18 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_18 <= _GEN_1194;
        end else begin
          predictor_18 <= _GEN_1322;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_18 <= _GEN_1834;
      end else begin
        predictor_18 <= _GEN_2858;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_19 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_19 <= _GEN_1195;
        end else begin
          predictor_19 <= _GEN_1323;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_19 <= _GEN_1835;
      end else begin
        predictor_19 <= _GEN_2859;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_20 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_20 <= _GEN_1196;
        end else begin
          predictor_20 <= _GEN_1324;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_20 <= _GEN_1836;
      end else begin
        predictor_20 <= _GEN_2860;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_21 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_21 <= _GEN_1197;
        end else begin
          predictor_21 <= _GEN_1325;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_21 <= _GEN_1837;
      end else begin
        predictor_21 <= _GEN_2861;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_22 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_22 <= _GEN_1198;
        end else begin
          predictor_22 <= _GEN_1326;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_22 <= _GEN_1838;
      end else begin
        predictor_22 <= _GEN_2862;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_23 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_23 <= _GEN_1199;
        end else begin
          predictor_23 <= _GEN_1327;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_23 <= _GEN_1839;
      end else begin
        predictor_23 <= _GEN_2863;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_24 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_24 <= _GEN_1200;
        end else begin
          predictor_24 <= _GEN_1328;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_24 <= _GEN_1840;
      end else begin
        predictor_24 <= _GEN_2864;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_25 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_25 <= _GEN_1201;
        end else begin
          predictor_25 <= _GEN_1329;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_25 <= _GEN_1841;
      end else begin
        predictor_25 <= _GEN_2865;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_26 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_26 <= _GEN_1202;
        end else begin
          predictor_26 <= _GEN_1330;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_26 <= _GEN_1842;
      end else begin
        predictor_26 <= _GEN_2866;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_27 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_27 <= _GEN_1203;
        end else begin
          predictor_27 <= _GEN_1331;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_27 <= _GEN_1843;
      end else begin
        predictor_27 <= _GEN_2867;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_28 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_28 <= _GEN_1204;
        end else begin
          predictor_28 <= _GEN_1332;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_28 <= _GEN_1844;
      end else begin
        predictor_28 <= _GEN_2868;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_29 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_29 <= _GEN_1205;
        end else begin
          predictor_29 <= _GEN_1333;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_29 <= _GEN_1845;
      end else begin
        predictor_29 <= _GEN_2869;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_30 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_30 <= _GEN_1206;
        end else begin
          predictor_30 <= _GEN_1334;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_30 <= _GEN_1846;
      end else begin
        predictor_30 <= _GEN_2870;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_31 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_31 <= _GEN_1207;
        end else begin
          predictor_31 <= _GEN_1335;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_31 <= _GEN_1847;
      end else begin
        predictor_31 <= _GEN_2871;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_32 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_32 <= _GEN_1208;
        end else begin
          predictor_32 <= _GEN_1336;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_32 <= _GEN_1848;
      end else begin
        predictor_32 <= _GEN_2872;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_33 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_33 <= _GEN_1209;
        end else begin
          predictor_33 <= _GEN_1337;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_33 <= _GEN_1849;
      end else begin
        predictor_33 <= _GEN_2873;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_34 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_34 <= _GEN_1210;
        end else begin
          predictor_34 <= _GEN_1338;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_34 <= _GEN_1850;
      end else begin
        predictor_34 <= _GEN_2874;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_35 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_35 <= _GEN_1211;
        end else begin
          predictor_35 <= _GEN_1339;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_35 <= _GEN_1851;
      end else begin
        predictor_35 <= _GEN_2875;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_36 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_36 <= _GEN_1212;
        end else begin
          predictor_36 <= _GEN_1340;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_36 <= _GEN_1852;
      end else begin
        predictor_36 <= _GEN_2876;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_37 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_37 <= _GEN_1213;
        end else begin
          predictor_37 <= _GEN_1341;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_37 <= _GEN_1853;
      end else begin
        predictor_37 <= _GEN_2877;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_38 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_38 <= _GEN_1214;
        end else begin
          predictor_38 <= _GEN_1342;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_38 <= _GEN_1854;
      end else begin
        predictor_38 <= _GEN_2878;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_39 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_39 <= _GEN_1215;
        end else begin
          predictor_39 <= _GEN_1343;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_39 <= _GEN_1855;
      end else begin
        predictor_39 <= _GEN_2879;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_40 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_40 <= _GEN_1216;
        end else begin
          predictor_40 <= _GEN_1344;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_40 <= _GEN_1856;
      end else begin
        predictor_40 <= _GEN_2880;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_41 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_41 <= _GEN_1217;
        end else begin
          predictor_41 <= _GEN_1345;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_41 <= _GEN_1857;
      end else begin
        predictor_41 <= _GEN_2881;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_42 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_42 <= _GEN_1218;
        end else begin
          predictor_42 <= _GEN_1346;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_42 <= _GEN_1858;
      end else begin
        predictor_42 <= _GEN_2882;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_43 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_43 <= _GEN_1219;
        end else begin
          predictor_43 <= _GEN_1347;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_43 <= _GEN_1859;
      end else begin
        predictor_43 <= _GEN_2883;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_44 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_44 <= _GEN_1220;
        end else begin
          predictor_44 <= _GEN_1348;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_44 <= _GEN_1860;
      end else begin
        predictor_44 <= _GEN_2884;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_45 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_45 <= _GEN_1221;
        end else begin
          predictor_45 <= _GEN_1349;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_45 <= _GEN_1861;
      end else begin
        predictor_45 <= _GEN_2885;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_46 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_46 <= _GEN_1222;
        end else begin
          predictor_46 <= _GEN_1350;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_46 <= _GEN_1862;
      end else begin
        predictor_46 <= _GEN_2886;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_47 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_47 <= _GEN_1223;
        end else begin
          predictor_47 <= _GEN_1351;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_47 <= _GEN_1863;
      end else begin
        predictor_47 <= _GEN_2887;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_48 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_48 <= _GEN_1224;
        end else begin
          predictor_48 <= _GEN_1352;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_48 <= _GEN_1864;
      end else begin
        predictor_48 <= _GEN_2888;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_49 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_49 <= _GEN_1225;
        end else begin
          predictor_49 <= _GEN_1353;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_49 <= _GEN_1865;
      end else begin
        predictor_49 <= _GEN_2889;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_50 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_50 <= _GEN_1226;
        end else begin
          predictor_50 <= _GEN_1354;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_50 <= _GEN_1866;
      end else begin
        predictor_50 <= _GEN_2890;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_51 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_51 <= _GEN_1227;
        end else begin
          predictor_51 <= _GEN_1355;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_51 <= _GEN_1867;
      end else begin
        predictor_51 <= _GEN_2891;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_52 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_52 <= _GEN_1228;
        end else begin
          predictor_52 <= _GEN_1356;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_52 <= _GEN_1868;
      end else begin
        predictor_52 <= _GEN_2892;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_53 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_53 <= _GEN_1229;
        end else begin
          predictor_53 <= _GEN_1357;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_53 <= _GEN_1869;
      end else begin
        predictor_53 <= _GEN_2893;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_54 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_54 <= _GEN_1230;
        end else begin
          predictor_54 <= _GEN_1358;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_54 <= _GEN_1870;
      end else begin
        predictor_54 <= _GEN_2894;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_55 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_55 <= _GEN_1231;
        end else begin
          predictor_55 <= _GEN_1359;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_55 <= _GEN_1871;
      end else begin
        predictor_55 <= _GEN_2895;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_56 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_56 <= _GEN_1232;
        end else begin
          predictor_56 <= _GEN_1360;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_56 <= _GEN_1872;
      end else begin
        predictor_56 <= _GEN_2896;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_57 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_57 <= _GEN_1233;
        end else begin
          predictor_57 <= _GEN_1361;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_57 <= _GEN_1873;
      end else begin
        predictor_57 <= _GEN_2897;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_58 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_58 <= _GEN_1234;
        end else begin
          predictor_58 <= _GEN_1362;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_58 <= _GEN_1874;
      end else begin
        predictor_58 <= _GEN_2898;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_59 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_59 <= _GEN_1235;
        end else begin
          predictor_59 <= _GEN_1363;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_59 <= _GEN_1875;
      end else begin
        predictor_59 <= _GEN_2899;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_60 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_60 <= _GEN_1236;
        end else begin
          predictor_60 <= _GEN_1364;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_60 <= _GEN_1876;
      end else begin
        predictor_60 <= _GEN_2900;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_61 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_61 <= _GEN_1237;
        end else begin
          predictor_61 <= _GEN_1365;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_61 <= _GEN_1877;
      end else begin
        predictor_61 <= _GEN_2901;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_62 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_62 <= _GEN_1238;
        end else begin
          predictor_62 <= _GEN_1366;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_62 <= _GEN_1878;
      end else begin
        predictor_62 <= _GEN_2902;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_63 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_63 <= _GEN_1239;
        end else begin
          predictor_63 <= _GEN_1367;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_63 <= _GEN_1879;
      end else begin
        predictor_63 <= _GEN_2903;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_64 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_64 <= _GEN_1240;
        end else begin
          predictor_64 <= _GEN_1368;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_64 <= _GEN_1880;
      end else begin
        predictor_64 <= _GEN_2904;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_65 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_65 <= _GEN_1241;
        end else begin
          predictor_65 <= _GEN_1369;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_65 <= _GEN_1881;
      end else begin
        predictor_65 <= _GEN_2905;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_66 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_66 <= _GEN_1242;
        end else begin
          predictor_66 <= _GEN_1370;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_66 <= _GEN_1882;
      end else begin
        predictor_66 <= _GEN_2906;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_67 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_67 <= _GEN_1243;
        end else begin
          predictor_67 <= _GEN_1371;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_67 <= _GEN_1883;
      end else begin
        predictor_67 <= _GEN_2907;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_68 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_68 <= _GEN_1244;
        end else begin
          predictor_68 <= _GEN_1372;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_68 <= _GEN_1884;
      end else begin
        predictor_68 <= _GEN_2908;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_69 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_69 <= _GEN_1245;
        end else begin
          predictor_69 <= _GEN_1373;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_69 <= _GEN_1885;
      end else begin
        predictor_69 <= _GEN_2909;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_70 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_70 <= _GEN_1246;
        end else begin
          predictor_70 <= _GEN_1374;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_70 <= _GEN_1886;
      end else begin
        predictor_70 <= _GEN_2910;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_71 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_71 <= _GEN_1247;
        end else begin
          predictor_71 <= _GEN_1375;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_71 <= _GEN_1887;
      end else begin
        predictor_71 <= _GEN_2911;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_72 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_72 <= _GEN_1248;
        end else begin
          predictor_72 <= _GEN_1376;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_72 <= _GEN_1888;
      end else begin
        predictor_72 <= _GEN_2912;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_73 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_73 <= _GEN_1249;
        end else begin
          predictor_73 <= _GEN_1377;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_73 <= _GEN_1889;
      end else begin
        predictor_73 <= _GEN_2913;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_74 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_74 <= _GEN_1250;
        end else begin
          predictor_74 <= _GEN_1378;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_74 <= _GEN_1890;
      end else begin
        predictor_74 <= _GEN_2914;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_75 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_75 <= _GEN_1251;
        end else begin
          predictor_75 <= _GEN_1379;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_75 <= _GEN_1891;
      end else begin
        predictor_75 <= _GEN_2915;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_76 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_76 <= _GEN_1252;
        end else begin
          predictor_76 <= _GEN_1380;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_76 <= _GEN_1892;
      end else begin
        predictor_76 <= _GEN_2916;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_77 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_77 <= _GEN_1253;
        end else begin
          predictor_77 <= _GEN_1381;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_77 <= _GEN_1893;
      end else begin
        predictor_77 <= _GEN_2917;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_78 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_78 <= _GEN_1254;
        end else begin
          predictor_78 <= _GEN_1382;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_78 <= _GEN_1894;
      end else begin
        predictor_78 <= _GEN_2918;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_79 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_79 <= _GEN_1255;
        end else begin
          predictor_79 <= _GEN_1383;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_79 <= _GEN_1895;
      end else begin
        predictor_79 <= _GEN_2919;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_80 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_80 <= _GEN_1256;
        end else begin
          predictor_80 <= _GEN_1384;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_80 <= _GEN_1896;
      end else begin
        predictor_80 <= _GEN_2920;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_81 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_81 <= _GEN_1257;
        end else begin
          predictor_81 <= _GEN_1385;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_81 <= _GEN_1897;
      end else begin
        predictor_81 <= _GEN_2921;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_82 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_82 <= _GEN_1258;
        end else begin
          predictor_82 <= _GEN_1386;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_82 <= _GEN_1898;
      end else begin
        predictor_82 <= _GEN_2922;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_83 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_83 <= _GEN_1259;
        end else begin
          predictor_83 <= _GEN_1387;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_83 <= _GEN_1899;
      end else begin
        predictor_83 <= _GEN_2923;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_84 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_84 <= _GEN_1260;
        end else begin
          predictor_84 <= _GEN_1388;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_84 <= _GEN_1900;
      end else begin
        predictor_84 <= _GEN_2924;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_85 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_85 <= _GEN_1261;
        end else begin
          predictor_85 <= _GEN_1389;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_85 <= _GEN_1901;
      end else begin
        predictor_85 <= _GEN_2925;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_86 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_86 <= _GEN_1262;
        end else begin
          predictor_86 <= _GEN_1390;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_86 <= _GEN_1902;
      end else begin
        predictor_86 <= _GEN_2926;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_87 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_87 <= _GEN_1263;
        end else begin
          predictor_87 <= _GEN_1391;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_87 <= _GEN_1903;
      end else begin
        predictor_87 <= _GEN_2927;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_88 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_88 <= _GEN_1264;
        end else begin
          predictor_88 <= _GEN_1392;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_88 <= _GEN_1904;
      end else begin
        predictor_88 <= _GEN_2928;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_89 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_89 <= _GEN_1265;
        end else begin
          predictor_89 <= _GEN_1393;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_89 <= _GEN_1905;
      end else begin
        predictor_89 <= _GEN_2929;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_90 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_90 <= _GEN_1266;
        end else begin
          predictor_90 <= _GEN_1394;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_90 <= _GEN_1906;
      end else begin
        predictor_90 <= _GEN_2930;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_91 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_91 <= _GEN_1267;
        end else begin
          predictor_91 <= _GEN_1395;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_91 <= _GEN_1907;
      end else begin
        predictor_91 <= _GEN_2931;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_92 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_92 <= _GEN_1268;
        end else begin
          predictor_92 <= _GEN_1396;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_92 <= _GEN_1908;
      end else begin
        predictor_92 <= _GEN_2932;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_93 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_93 <= _GEN_1269;
        end else begin
          predictor_93 <= _GEN_1397;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_93 <= _GEN_1909;
      end else begin
        predictor_93 <= _GEN_2933;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_94 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_94 <= _GEN_1270;
        end else begin
          predictor_94 <= _GEN_1398;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_94 <= _GEN_1910;
      end else begin
        predictor_94 <= _GEN_2934;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_95 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_95 <= _GEN_1271;
        end else begin
          predictor_95 <= _GEN_1399;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_95 <= _GEN_1911;
      end else begin
        predictor_95 <= _GEN_2935;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_96 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_96 <= _GEN_1272;
        end else begin
          predictor_96 <= _GEN_1400;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_96 <= _GEN_1912;
      end else begin
        predictor_96 <= _GEN_2936;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_97 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_97 <= _GEN_1273;
        end else begin
          predictor_97 <= _GEN_1401;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_97 <= _GEN_1913;
      end else begin
        predictor_97 <= _GEN_2937;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_98 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_98 <= _GEN_1274;
        end else begin
          predictor_98 <= _GEN_1402;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_98 <= _GEN_1914;
      end else begin
        predictor_98 <= _GEN_2938;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_99 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_99 <= _GEN_1275;
        end else begin
          predictor_99 <= _GEN_1403;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_99 <= _GEN_1915;
      end else begin
        predictor_99 <= _GEN_2939;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_100 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_100 <= _GEN_1276;
        end else begin
          predictor_100 <= _GEN_1404;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_100 <= _GEN_1916;
      end else begin
        predictor_100 <= _GEN_2940;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_101 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_101 <= _GEN_1277;
        end else begin
          predictor_101 <= _GEN_1405;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_101 <= _GEN_1917;
      end else begin
        predictor_101 <= _GEN_2941;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_102 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_102 <= _GEN_1278;
        end else begin
          predictor_102 <= _GEN_1406;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_102 <= _GEN_1918;
      end else begin
        predictor_102 <= _GEN_2942;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_103 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_103 <= _GEN_1279;
        end else begin
          predictor_103 <= _GEN_1407;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_103 <= _GEN_1919;
      end else begin
        predictor_103 <= _GEN_2943;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_104 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_104 <= _GEN_1280;
        end else begin
          predictor_104 <= _GEN_1408;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_104 <= _GEN_1920;
      end else begin
        predictor_104 <= _GEN_2944;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_105 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_105 <= _GEN_1281;
        end else begin
          predictor_105 <= _GEN_1409;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_105 <= _GEN_1921;
      end else begin
        predictor_105 <= _GEN_2945;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_106 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_106 <= _GEN_1282;
        end else begin
          predictor_106 <= _GEN_1410;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_106 <= _GEN_1922;
      end else begin
        predictor_106 <= _GEN_2946;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_107 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_107 <= _GEN_1283;
        end else begin
          predictor_107 <= _GEN_1411;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_107 <= _GEN_1923;
      end else begin
        predictor_107 <= _GEN_2947;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_108 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_108 <= _GEN_1284;
        end else begin
          predictor_108 <= _GEN_1412;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_108 <= _GEN_1924;
      end else begin
        predictor_108 <= _GEN_2948;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_109 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_109 <= _GEN_1285;
        end else begin
          predictor_109 <= _GEN_1413;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_109 <= _GEN_1925;
      end else begin
        predictor_109 <= _GEN_2949;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_110 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_110 <= _GEN_1286;
        end else begin
          predictor_110 <= _GEN_1414;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_110 <= _GEN_1926;
      end else begin
        predictor_110 <= _GEN_2950;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_111 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_111 <= _GEN_1287;
        end else begin
          predictor_111 <= _GEN_1415;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_111 <= _GEN_1927;
      end else begin
        predictor_111 <= _GEN_2951;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_112 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_112 <= _GEN_1288;
        end else begin
          predictor_112 <= _GEN_1416;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_112 <= _GEN_1928;
      end else begin
        predictor_112 <= _GEN_2952;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_113 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_113 <= _GEN_1289;
        end else begin
          predictor_113 <= _GEN_1417;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_113 <= _GEN_1929;
      end else begin
        predictor_113 <= _GEN_2953;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_114 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_114 <= _GEN_1290;
        end else begin
          predictor_114 <= _GEN_1418;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_114 <= _GEN_1930;
      end else begin
        predictor_114 <= _GEN_2954;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_115 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_115 <= _GEN_1291;
        end else begin
          predictor_115 <= _GEN_1419;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_115 <= _GEN_1931;
      end else begin
        predictor_115 <= _GEN_2955;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_116 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_116 <= _GEN_1292;
        end else begin
          predictor_116 <= _GEN_1420;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_116 <= _GEN_1932;
      end else begin
        predictor_116 <= _GEN_2956;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_117 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_117 <= _GEN_1293;
        end else begin
          predictor_117 <= _GEN_1421;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_117 <= _GEN_1933;
      end else begin
        predictor_117 <= _GEN_2957;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_118 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_118 <= _GEN_1294;
        end else begin
          predictor_118 <= _GEN_1422;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_118 <= _GEN_1934;
      end else begin
        predictor_118 <= _GEN_2958;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_119 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_119 <= _GEN_1295;
        end else begin
          predictor_119 <= _GEN_1423;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_119 <= _GEN_1935;
      end else begin
        predictor_119 <= _GEN_2959;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_120 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_120 <= _GEN_1296;
        end else begin
          predictor_120 <= _GEN_1424;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_120 <= _GEN_1936;
      end else begin
        predictor_120 <= _GEN_2960;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_121 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_121 <= _GEN_1297;
        end else begin
          predictor_121 <= _GEN_1425;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_121 <= _GEN_1937;
      end else begin
        predictor_121 <= _GEN_2961;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_122 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_122 <= _GEN_1298;
        end else begin
          predictor_122 <= _GEN_1426;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_122 <= _GEN_1938;
      end else begin
        predictor_122 <= _GEN_2962;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_123 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_123 <= _GEN_1299;
        end else begin
          predictor_123 <= _GEN_1427;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_123 <= _GEN_1939;
      end else begin
        predictor_123 <= _GEN_2963;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_124 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_124 <= _GEN_1300;
        end else begin
          predictor_124 <= _GEN_1428;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_124 <= _GEN_1940;
      end else begin
        predictor_124 <= _GEN_2964;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_125 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_125 <= _GEN_1301;
        end else begin
          predictor_125 <= _GEN_1429;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_125 <= _GEN_1941;
      end else begin
        predictor_125 <= _GEN_2965;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_126 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_126 <= _GEN_1302;
        end else begin
          predictor_126 <= _GEN_1430;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_126 <= _GEN_1942;
      end else begin
        predictor_126 <= _GEN_2966;
      end
    end
    if (reset) begin // @[Bpu.scala 74:31]
      predictor_127 <= 2'h2; // @[Bpu.scala 74:31]
    end else if (io_branch_info_i_valid & io_branch_info_i_bits_is_branch) begin // @[Bpu.scala 127:67]
      if (_T_3) begin // @[Conditional.scala 40:58]
        if (io_branch_info_i_bits_is_taken) begin // @[Bpu.scala 130:46]
          predictor_127 <= _GEN_1303;
        end else begin
          predictor_127 <= _GEN_1431;
        end
      end else if (_T_4) begin // @[Conditional.scala 39:67]
        predictor_127 <= _GEN_1943;
      end else begin
        predictor_127 <= _GEN_2967;
      end
    end
    if (reset) begin // @[Bpu.scala 196:23]
      bpu_inst_packet_o_data_0 <= 32'h0; // @[Bpu.scala 17:18]
    end else if (io_need_flush) begin // @[Bpu.scala 191:22]
      bpu_inst_packet_o_data_0 <= 32'h0; // @[Bpu.scala 17:18]
    end else if (io_bpu_inst_packet_o_ready) begin // @[Bpu.scala 168:35]
      bpu_inst_packet_o_data_0 <= io_inst_packet_i_bits_data_0; // @[Bpu.scala 172:28]
    end
    if (reset) begin // @[Bpu.scala 196:23]
      bpu_inst_packet_o_data_1 <= 32'h0; // @[Bpu.scala 17:18]
    end else if (io_need_flush) begin // @[Bpu.scala 191:22]
      bpu_inst_packet_o_data_1 <= 32'h0; // @[Bpu.scala 17:18]
    end else if (io_bpu_inst_packet_o_ready) begin // @[Bpu.scala 168:35]
      bpu_inst_packet_o_data_1 <= io_inst_packet_i_bits_data_1; // @[Bpu.scala 172:28]
    end
    if (reset) begin // @[Bpu.scala 196:23]
      bpu_inst_packet_o_data_2 <= 32'h0; // @[Bpu.scala 17:18]
    end else if (io_need_flush) begin // @[Bpu.scala 191:22]
      bpu_inst_packet_o_data_2 <= 32'h0; // @[Bpu.scala 17:18]
    end else if (io_bpu_inst_packet_o_ready) begin // @[Bpu.scala 168:35]
      bpu_inst_packet_o_data_2 <= io_inst_packet_i_bits_data_2; // @[Bpu.scala 172:28]
    end
    if (reset) begin // @[Bpu.scala 196:23]
      bpu_inst_packet_o_data_3 <= 32'h0; // @[Bpu.scala 17:18]
    end else if (io_need_flush) begin // @[Bpu.scala 191:22]
      bpu_inst_packet_o_data_3 <= 32'h0; // @[Bpu.scala 17:18]
    end else if (io_bpu_inst_packet_o_ready) begin // @[Bpu.scala 168:35]
      bpu_inst_packet_o_data_3 <= io_inst_packet_i_bits_data_3; // @[Bpu.scala 172:28]
    end
    if (reset) begin // @[Bpu.scala 196:23]
      bpu_inst_packet_o_data_4 <= 32'h0; // @[Bpu.scala 17:18]
    end else if (io_need_flush) begin // @[Bpu.scala 191:22]
      bpu_inst_packet_o_data_4 <= 32'h0; // @[Bpu.scala 17:18]
    end else if (io_bpu_inst_packet_o_ready) begin // @[Bpu.scala 168:35]
      bpu_inst_packet_o_data_4 <= io_inst_packet_i_bits_data_4; // @[Bpu.scala 172:28]
    end
    if (reset) begin // @[Bpu.scala 196:23]
      bpu_inst_packet_o_data_5 <= 32'h0; // @[Bpu.scala 17:18]
    end else if (io_need_flush) begin // @[Bpu.scala 191:22]
      bpu_inst_packet_o_data_5 <= 32'h0; // @[Bpu.scala 17:18]
    end else if (io_bpu_inst_packet_o_ready) begin // @[Bpu.scala 168:35]
      bpu_inst_packet_o_data_5 <= io_inst_packet_i_bits_data_5; // @[Bpu.scala 172:28]
    end
    if (reset) begin // @[Bpu.scala 196:23]
      bpu_inst_packet_o_data_6 <= 32'h0; // @[Bpu.scala 17:18]
    end else if (io_need_flush) begin // @[Bpu.scala 191:22]
      bpu_inst_packet_o_data_6 <= 32'h0; // @[Bpu.scala 17:18]
    end else if (io_bpu_inst_packet_o_ready) begin // @[Bpu.scala 168:35]
      bpu_inst_packet_o_data_6 <= io_inst_packet_i_bits_data_6; // @[Bpu.scala 172:28]
    end
    if (reset) begin // @[Bpu.scala 196:23]
      bpu_inst_packet_o_data_7 <= 32'h0; // @[Bpu.scala 17:18]
    end else if (io_need_flush) begin // @[Bpu.scala 191:22]
      bpu_inst_packet_o_data_7 <= 32'h0; // @[Bpu.scala 17:18]
    end else if (io_bpu_inst_packet_o_ready) begin // @[Bpu.scala 168:35]
      bpu_inst_packet_o_data_7 <= io_inst_packet_i_bits_data_7; // @[Bpu.scala 172:28]
    end
    if (reset) begin // @[Bpu.scala 196:23]
      bpu_inst_packet_o_addr <= 32'h0; // @[Bpu.scala 18:18]
    end else if (io_need_flush) begin // @[Bpu.scala 191:22]
      bpu_inst_packet_o_addr <= 32'h0; // @[Bpu.scala 18:18]
    end else if (io_bpu_inst_packet_o_ready) begin // @[Bpu.scala 168:35]
      bpu_inst_packet_o_addr <= io_inst_packet_i_bits_addr; // @[Bpu.scala 171:28]
    end
    if (reset) begin // @[Bpu.scala 196:23]
      bpu_inst_packet_o_gh_backup <= 4'h0; // @[Bpu.scala 19:18]
    end else if (io_need_flush) begin // @[Bpu.scala 191:22]
      bpu_inst_packet_o_gh_backup <= 4'h0; // @[Bpu.scala 19:18]
    end else if (io_bpu_inst_packet_o_ready) begin // @[Bpu.scala 168:35]
      bpu_inst_packet_o_gh_backup <= global_history; // @[Bpu.scala 176:33]
    end
    if (reset) begin // @[Bpu.scala 196:23]
      bpu_inst_packet_o_valid_mask_0 <= 1'h0; // @[Bpu.scala 20:18]
    end else if (io_need_flush) begin // @[Bpu.scala 191:22]
      bpu_inst_packet_o_valid_mask_0 <= 1'h0; // @[Bpu.scala 20:18]
    end else if (io_bpu_inst_packet_o_ready) begin // @[Bpu.scala 168:35]
      if (~take_delay & is_taken) begin // @[Bpu.scala 121:33]
        bpu_inst_packet_o_valid_mask_0 <= _GEN_1032;
      end else begin
        bpu_inst_packet_o_valid_mask_0 <= (inst_mask_0 | (inst_mask_1 | (inst_mask_2 | (inst_mask_3 | (inst_mask_4 | (
          inst_mask_5 | (inst_mask_6 | (inst_mask_7 | ~is_taken)))))))) & fetched_mask_0; // @[Bpu.scala 119:27]
      end
    end
    if (reset) begin // @[Bpu.scala 196:23]
      bpu_inst_packet_o_valid_mask_1 <= 1'h0; // @[Bpu.scala 20:18]
    end else if (io_need_flush) begin // @[Bpu.scala 191:22]
      bpu_inst_packet_o_valid_mask_1 <= 1'h0; // @[Bpu.scala 20:18]
    end else if (io_bpu_inst_packet_o_ready) begin // @[Bpu.scala 168:35]
      if (~take_delay & is_taken) begin // @[Bpu.scala 121:33]
        bpu_inst_packet_o_valid_mask_1 <= _GEN_1033;
      end else begin
        bpu_inst_packet_o_valid_mask_1 <= (inst_mask_1 | (inst_mask_2 | (inst_mask_3 | (inst_mask_4 | (inst_mask_5 | (
          inst_mask_6 | (inst_mask_7 | ~is_taken))))))) & fetched_mask_1; // @[Bpu.scala 119:27]
      end
    end
    if (reset) begin // @[Bpu.scala 196:23]
      bpu_inst_packet_o_valid_mask_2 <= 1'h0; // @[Bpu.scala 20:18]
    end else if (io_need_flush) begin // @[Bpu.scala 191:22]
      bpu_inst_packet_o_valid_mask_2 <= 1'h0; // @[Bpu.scala 20:18]
    end else if (io_bpu_inst_packet_o_ready) begin // @[Bpu.scala 168:35]
      if (~take_delay & is_taken) begin // @[Bpu.scala 121:33]
        bpu_inst_packet_o_valid_mask_2 <= _GEN_1034;
      end else begin
        bpu_inst_packet_o_valid_mask_2 <= (inst_mask_2 | (inst_mask_3 | (inst_mask_4 | (inst_mask_5 | (inst_mask_6 | (
          inst_mask_7 | ~is_taken)))))) & fetched_mask_2; // @[Bpu.scala 119:27]
      end
    end
    if (reset) begin // @[Bpu.scala 196:23]
      bpu_inst_packet_o_valid_mask_3 <= 1'h0; // @[Bpu.scala 20:18]
    end else if (io_need_flush) begin // @[Bpu.scala 191:22]
      bpu_inst_packet_o_valid_mask_3 <= 1'h0; // @[Bpu.scala 20:18]
    end else if (io_bpu_inst_packet_o_ready) begin // @[Bpu.scala 168:35]
      if (~take_delay & is_taken) begin // @[Bpu.scala 121:33]
        bpu_inst_packet_o_valid_mask_3 <= _GEN_1035;
      end else begin
        bpu_inst_packet_o_valid_mask_3 <= (inst_mask_3 | (inst_mask_4 | (inst_mask_5 | (inst_mask_6 | (inst_mask_7 | ~
          is_taken))))) & fetched_mask_3; // @[Bpu.scala 119:27]
      end
    end
    if (reset) begin // @[Bpu.scala 196:23]
      bpu_inst_packet_o_valid_mask_4 <= 1'h0; // @[Bpu.scala 20:18]
    end else if (io_need_flush) begin // @[Bpu.scala 191:22]
      bpu_inst_packet_o_valid_mask_4 <= 1'h0; // @[Bpu.scala 20:18]
    end else if (io_bpu_inst_packet_o_ready) begin // @[Bpu.scala 168:35]
      if (~take_delay & is_taken) begin // @[Bpu.scala 121:33]
        bpu_inst_packet_o_valid_mask_4 <= _GEN_1036;
      end else begin
        bpu_inst_packet_o_valid_mask_4 <= (inst_mask_4 | (inst_mask_5 | (inst_mask_6 | (inst_mask_7 | ~is_taken)))) &
          fetched_mask_4; // @[Bpu.scala 119:27]
      end
    end
    if (reset) begin // @[Bpu.scala 196:23]
      bpu_inst_packet_o_valid_mask_5 <= 1'h0; // @[Bpu.scala 20:18]
    end else if (io_need_flush) begin // @[Bpu.scala 191:22]
      bpu_inst_packet_o_valid_mask_5 <= 1'h0; // @[Bpu.scala 20:18]
    end else if (io_bpu_inst_packet_o_ready) begin // @[Bpu.scala 168:35]
      if (~take_delay & is_taken) begin // @[Bpu.scala 121:33]
        bpu_inst_packet_o_valid_mask_5 <= _GEN_1037;
      end else begin
        bpu_inst_packet_o_valid_mask_5 <= (inst_mask_5 | (inst_mask_6 | (inst_mask_7 | ~is_taken))) & fetched_mask_5; // @[Bpu.scala 119:27]
      end
    end
    if (reset) begin // @[Bpu.scala 196:23]
      bpu_inst_packet_o_valid_mask_6 <= 1'h0; // @[Bpu.scala 20:18]
    end else if (io_need_flush) begin // @[Bpu.scala 191:22]
      bpu_inst_packet_o_valid_mask_6 <= 1'h0; // @[Bpu.scala 20:18]
    end else if (io_bpu_inst_packet_o_ready) begin // @[Bpu.scala 168:35]
      if (~take_delay & is_taken) begin // @[Bpu.scala 121:33]
        bpu_inst_packet_o_valid_mask_6 <= _GEN_1038;
      end else begin
        bpu_inst_packet_o_valid_mask_6 <= (inst_mask_6 | (inst_mask_7 | ~is_taken)) & fetched_mask_6; // @[Bpu.scala 119:27]
      end
    end
    if (reset) begin // @[Bpu.scala 196:23]
      bpu_inst_packet_o_valid_mask_7 <= 1'h0; // @[Bpu.scala 20:18]
    end else if (io_need_flush) begin // @[Bpu.scala 191:22]
      bpu_inst_packet_o_valid_mask_7 <= 1'h0; // @[Bpu.scala 20:18]
    end else if (io_bpu_inst_packet_o_ready) begin // @[Bpu.scala 168:35]
      if (~take_delay & is_taken) begin // @[Bpu.scala 121:33]
        bpu_inst_packet_o_valid_mask_7 <= _GEN_1039;
      end else begin
        bpu_inst_packet_o_valid_mask_7 <= (inst_mask_7 | ~is_taken) & fetched_mask_7; // @[Bpu.scala 119:27]
      end
    end
    if (reset) begin // @[Bpu.scala 196:23]
      bpu_inst_packet_o_predict_mask_0 <= 1'h0; // @[Bpu.scala 23:19]
    end else if (io_need_flush) begin // @[Bpu.scala 191:22]
      bpu_inst_packet_o_predict_mask_0 <= 1'h0; // @[Bpu.scala 23:19]
    end else if (io_bpu_inst_packet_o_ready) begin // @[Bpu.scala 168:35]
      bpu_inst_packet_o_predict_mask_0 <= predict_branch_0; // @[Bpu.scala 174:36]
    end
    if (reset) begin // @[Bpu.scala 196:23]
      bpu_inst_packet_o_predict_mask_1 <= 1'h0; // @[Bpu.scala 23:19]
    end else if (io_need_flush) begin // @[Bpu.scala 191:22]
      bpu_inst_packet_o_predict_mask_1 <= 1'h0; // @[Bpu.scala 23:19]
    end else if (io_bpu_inst_packet_o_ready) begin // @[Bpu.scala 168:35]
      bpu_inst_packet_o_predict_mask_1 <= predict_branch_1; // @[Bpu.scala 174:36]
    end
    if (reset) begin // @[Bpu.scala 196:23]
      bpu_inst_packet_o_predict_mask_2 <= 1'h0; // @[Bpu.scala 23:19]
    end else if (io_need_flush) begin // @[Bpu.scala 191:22]
      bpu_inst_packet_o_predict_mask_2 <= 1'h0; // @[Bpu.scala 23:19]
    end else if (io_bpu_inst_packet_o_ready) begin // @[Bpu.scala 168:35]
      bpu_inst_packet_o_predict_mask_2 <= predict_branch_2; // @[Bpu.scala 174:36]
    end
    if (reset) begin // @[Bpu.scala 196:23]
      bpu_inst_packet_o_predict_mask_3 <= 1'h0; // @[Bpu.scala 23:19]
    end else if (io_need_flush) begin // @[Bpu.scala 191:22]
      bpu_inst_packet_o_predict_mask_3 <= 1'h0; // @[Bpu.scala 23:19]
    end else if (io_bpu_inst_packet_o_ready) begin // @[Bpu.scala 168:35]
      bpu_inst_packet_o_predict_mask_3 <= predict_branch_3; // @[Bpu.scala 174:36]
    end
    if (reset) begin // @[Bpu.scala 196:23]
      bpu_inst_packet_o_predict_mask_4 <= 1'h0; // @[Bpu.scala 23:19]
    end else if (io_need_flush) begin // @[Bpu.scala 191:22]
      bpu_inst_packet_o_predict_mask_4 <= 1'h0; // @[Bpu.scala 23:19]
    end else if (io_bpu_inst_packet_o_ready) begin // @[Bpu.scala 168:35]
      bpu_inst_packet_o_predict_mask_4 <= predict_branch_4; // @[Bpu.scala 174:36]
    end
    if (reset) begin // @[Bpu.scala 196:23]
      bpu_inst_packet_o_predict_mask_5 <= 1'h0; // @[Bpu.scala 23:19]
    end else if (io_need_flush) begin // @[Bpu.scala 191:22]
      bpu_inst_packet_o_predict_mask_5 <= 1'h0; // @[Bpu.scala 23:19]
    end else if (io_bpu_inst_packet_o_ready) begin // @[Bpu.scala 168:35]
      bpu_inst_packet_o_predict_mask_5 <= predict_branch_5; // @[Bpu.scala 174:36]
    end
    if (reset) begin // @[Bpu.scala 196:23]
      bpu_inst_packet_o_predict_mask_6 <= 1'h0; // @[Bpu.scala 23:19]
    end else if (io_need_flush) begin // @[Bpu.scala 191:22]
      bpu_inst_packet_o_predict_mask_6 <= 1'h0; // @[Bpu.scala 23:19]
    end else if (io_bpu_inst_packet_o_ready) begin // @[Bpu.scala 168:35]
      bpu_inst_packet_o_predict_mask_6 <= predict_branch_6; // @[Bpu.scala 174:36]
    end
    if (reset) begin // @[Bpu.scala 196:23]
      bpu_inst_packet_o_predict_mask_7 <= 1'h0; // @[Bpu.scala 23:19]
    end else if (io_need_flush) begin // @[Bpu.scala 191:22]
      bpu_inst_packet_o_predict_mask_7 <= 1'h0; // @[Bpu.scala 23:19]
    end else if (io_bpu_inst_packet_o_ready) begin // @[Bpu.scala 168:35]
      bpu_inst_packet_o_predict_mask_7 <= predict_branch_7; // @[Bpu.scala 174:36]
    end
    if (reset) begin // @[Bpu.scala 166:40]
      bpu_inst_packet_o_valid <= 1'h0; // @[Bpu.scala 166:40]
    end else if (io_need_flush) begin // @[Bpu.scala 191:22]
      bpu_inst_packet_o_valid <= 1'h0; // @[Bpu.scala 193:28]
    end else if (io_bpu_inst_packet_o_ready) begin // @[Bpu.scala 168:35]
      bpu_inst_packet_o_valid <= io_inst_packet_i_valid; // @[Bpu.scala 169:29]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  global_history = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  predictor_0 = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  predictor_1 = _RAND_2[1:0];
  _RAND_3 = {1{`RANDOM}};
  predictor_2 = _RAND_3[1:0];
  _RAND_4 = {1{`RANDOM}};
  predictor_3 = _RAND_4[1:0];
  _RAND_5 = {1{`RANDOM}};
  predictor_4 = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  predictor_5 = _RAND_6[1:0];
  _RAND_7 = {1{`RANDOM}};
  predictor_6 = _RAND_7[1:0];
  _RAND_8 = {1{`RANDOM}};
  predictor_7 = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  predictor_8 = _RAND_9[1:0];
  _RAND_10 = {1{`RANDOM}};
  predictor_9 = _RAND_10[1:0];
  _RAND_11 = {1{`RANDOM}};
  predictor_10 = _RAND_11[1:0];
  _RAND_12 = {1{`RANDOM}};
  predictor_11 = _RAND_12[1:0];
  _RAND_13 = {1{`RANDOM}};
  predictor_12 = _RAND_13[1:0];
  _RAND_14 = {1{`RANDOM}};
  predictor_13 = _RAND_14[1:0];
  _RAND_15 = {1{`RANDOM}};
  predictor_14 = _RAND_15[1:0];
  _RAND_16 = {1{`RANDOM}};
  predictor_15 = _RAND_16[1:0];
  _RAND_17 = {1{`RANDOM}};
  predictor_16 = _RAND_17[1:0];
  _RAND_18 = {1{`RANDOM}};
  predictor_17 = _RAND_18[1:0];
  _RAND_19 = {1{`RANDOM}};
  predictor_18 = _RAND_19[1:0];
  _RAND_20 = {1{`RANDOM}};
  predictor_19 = _RAND_20[1:0];
  _RAND_21 = {1{`RANDOM}};
  predictor_20 = _RAND_21[1:0];
  _RAND_22 = {1{`RANDOM}};
  predictor_21 = _RAND_22[1:0];
  _RAND_23 = {1{`RANDOM}};
  predictor_22 = _RAND_23[1:0];
  _RAND_24 = {1{`RANDOM}};
  predictor_23 = _RAND_24[1:0];
  _RAND_25 = {1{`RANDOM}};
  predictor_24 = _RAND_25[1:0];
  _RAND_26 = {1{`RANDOM}};
  predictor_25 = _RAND_26[1:0];
  _RAND_27 = {1{`RANDOM}};
  predictor_26 = _RAND_27[1:0];
  _RAND_28 = {1{`RANDOM}};
  predictor_27 = _RAND_28[1:0];
  _RAND_29 = {1{`RANDOM}};
  predictor_28 = _RAND_29[1:0];
  _RAND_30 = {1{`RANDOM}};
  predictor_29 = _RAND_30[1:0];
  _RAND_31 = {1{`RANDOM}};
  predictor_30 = _RAND_31[1:0];
  _RAND_32 = {1{`RANDOM}};
  predictor_31 = _RAND_32[1:0];
  _RAND_33 = {1{`RANDOM}};
  predictor_32 = _RAND_33[1:0];
  _RAND_34 = {1{`RANDOM}};
  predictor_33 = _RAND_34[1:0];
  _RAND_35 = {1{`RANDOM}};
  predictor_34 = _RAND_35[1:0];
  _RAND_36 = {1{`RANDOM}};
  predictor_35 = _RAND_36[1:0];
  _RAND_37 = {1{`RANDOM}};
  predictor_36 = _RAND_37[1:0];
  _RAND_38 = {1{`RANDOM}};
  predictor_37 = _RAND_38[1:0];
  _RAND_39 = {1{`RANDOM}};
  predictor_38 = _RAND_39[1:0];
  _RAND_40 = {1{`RANDOM}};
  predictor_39 = _RAND_40[1:0];
  _RAND_41 = {1{`RANDOM}};
  predictor_40 = _RAND_41[1:0];
  _RAND_42 = {1{`RANDOM}};
  predictor_41 = _RAND_42[1:0];
  _RAND_43 = {1{`RANDOM}};
  predictor_42 = _RAND_43[1:0];
  _RAND_44 = {1{`RANDOM}};
  predictor_43 = _RAND_44[1:0];
  _RAND_45 = {1{`RANDOM}};
  predictor_44 = _RAND_45[1:0];
  _RAND_46 = {1{`RANDOM}};
  predictor_45 = _RAND_46[1:0];
  _RAND_47 = {1{`RANDOM}};
  predictor_46 = _RAND_47[1:0];
  _RAND_48 = {1{`RANDOM}};
  predictor_47 = _RAND_48[1:0];
  _RAND_49 = {1{`RANDOM}};
  predictor_48 = _RAND_49[1:0];
  _RAND_50 = {1{`RANDOM}};
  predictor_49 = _RAND_50[1:0];
  _RAND_51 = {1{`RANDOM}};
  predictor_50 = _RAND_51[1:0];
  _RAND_52 = {1{`RANDOM}};
  predictor_51 = _RAND_52[1:0];
  _RAND_53 = {1{`RANDOM}};
  predictor_52 = _RAND_53[1:0];
  _RAND_54 = {1{`RANDOM}};
  predictor_53 = _RAND_54[1:0];
  _RAND_55 = {1{`RANDOM}};
  predictor_54 = _RAND_55[1:0];
  _RAND_56 = {1{`RANDOM}};
  predictor_55 = _RAND_56[1:0];
  _RAND_57 = {1{`RANDOM}};
  predictor_56 = _RAND_57[1:0];
  _RAND_58 = {1{`RANDOM}};
  predictor_57 = _RAND_58[1:0];
  _RAND_59 = {1{`RANDOM}};
  predictor_58 = _RAND_59[1:0];
  _RAND_60 = {1{`RANDOM}};
  predictor_59 = _RAND_60[1:0];
  _RAND_61 = {1{`RANDOM}};
  predictor_60 = _RAND_61[1:0];
  _RAND_62 = {1{`RANDOM}};
  predictor_61 = _RAND_62[1:0];
  _RAND_63 = {1{`RANDOM}};
  predictor_62 = _RAND_63[1:0];
  _RAND_64 = {1{`RANDOM}};
  predictor_63 = _RAND_64[1:0];
  _RAND_65 = {1{`RANDOM}};
  predictor_64 = _RAND_65[1:0];
  _RAND_66 = {1{`RANDOM}};
  predictor_65 = _RAND_66[1:0];
  _RAND_67 = {1{`RANDOM}};
  predictor_66 = _RAND_67[1:0];
  _RAND_68 = {1{`RANDOM}};
  predictor_67 = _RAND_68[1:0];
  _RAND_69 = {1{`RANDOM}};
  predictor_68 = _RAND_69[1:0];
  _RAND_70 = {1{`RANDOM}};
  predictor_69 = _RAND_70[1:0];
  _RAND_71 = {1{`RANDOM}};
  predictor_70 = _RAND_71[1:0];
  _RAND_72 = {1{`RANDOM}};
  predictor_71 = _RAND_72[1:0];
  _RAND_73 = {1{`RANDOM}};
  predictor_72 = _RAND_73[1:0];
  _RAND_74 = {1{`RANDOM}};
  predictor_73 = _RAND_74[1:0];
  _RAND_75 = {1{`RANDOM}};
  predictor_74 = _RAND_75[1:0];
  _RAND_76 = {1{`RANDOM}};
  predictor_75 = _RAND_76[1:0];
  _RAND_77 = {1{`RANDOM}};
  predictor_76 = _RAND_77[1:0];
  _RAND_78 = {1{`RANDOM}};
  predictor_77 = _RAND_78[1:0];
  _RAND_79 = {1{`RANDOM}};
  predictor_78 = _RAND_79[1:0];
  _RAND_80 = {1{`RANDOM}};
  predictor_79 = _RAND_80[1:0];
  _RAND_81 = {1{`RANDOM}};
  predictor_80 = _RAND_81[1:0];
  _RAND_82 = {1{`RANDOM}};
  predictor_81 = _RAND_82[1:0];
  _RAND_83 = {1{`RANDOM}};
  predictor_82 = _RAND_83[1:0];
  _RAND_84 = {1{`RANDOM}};
  predictor_83 = _RAND_84[1:0];
  _RAND_85 = {1{`RANDOM}};
  predictor_84 = _RAND_85[1:0];
  _RAND_86 = {1{`RANDOM}};
  predictor_85 = _RAND_86[1:0];
  _RAND_87 = {1{`RANDOM}};
  predictor_86 = _RAND_87[1:0];
  _RAND_88 = {1{`RANDOM}};
  predictor_87 = _RAND_88[1:0];
  _RAND_89 = {1{`RANDOM}};
  predictor_88 = _RAND_89[1:0];
  _RAND_90 = {1{`RANDOM}};
  predictor_89 = _RAND_90[1:0];
  _RAND_91 = {1{`RANDOM}};
  predictor_90 = _RAND_91[1:0];
  _RAND_92 = {1{`RANDOM}};
  predictor_91 = _RAND_92[1:0];
  _RAND_93 = {1{`RANDOM}};
  predictor_92 = _RAND_93[1:0];
  _RAND_94 = {1{`RANDOM}};
  predictor_93 = _RAND_94[1:0];
  _RAND_95 = {1{`RANDOM}};
  predictor_94 = _RAND_95[1:0];
  _RAND_96 = {1{`RANDOM}};
  predictor_95 = _RAND_96[1:0];
  _RAND_97 = {1{`RANDOM}};
  predictor_96 = _RAND_97[1:0];
  _RAND_98 = {1{`RANDOM}};
  predictor_97 = _RAND_98[1:0];
  _RAND_99 = {1{`RANDOM}};
  predictor_98 = _RAND_99[1:0];
  _RAND_100 = {1{`RANDOM}};
  predictor_99 = _RAND_100[1:0];
  _RAND_101 = {1{`RANDOM}};
  predictor_100 = _RAND_101[1:0];
  _RAND_102 = {1{`RANDOM}};
  predictor_101 = _RAND_102[1:0];
  _RAND_103 = {1{`RANDOM}};
  predictor_102 = _RAND_103[1:0];
  _RAND_104 = {1{`RANDOM}};
  predictor_103 = _RAND_104[1:0];
  _RAND_105 = {1{`RANDOM}};
  predictor_104 = _RAND_105[1:0];
  _RAND_106 = {1{`RANDOM}};
  predictor_105 = _RAND_106[1:0];
  _RAND_107 = {1{`RANDOM}};
  predictor_106 = _RAND_107[1:0];
  _RAND_108 = {1{`RANDOM}};
  predictor_107 = _RAND_108[1:0];
  _RAND_109 = {1{`RANDOM}};
  predictor_108 = _RAND_109[1:0];
  _RAND_110 = {1{`RANDOM}};
  predictor_109 = _RAND_110[1:0];
  _RAND_111 = {1{`RANDOM}};
  predictor_110 = _RAND_111[1:0];
  _RAND_112 = {1{`RANDOM}};
  predictor_111 = _RAND_112[1:0];
  _RAND_113 = {1{`RANDOM}};
  predictor_112 = _RAND_113[1:0];
  _RAND_114 = {1{`RANDOM}};
  predictor_113 = _RAND_114[1:0];
  _RAND_115 = {1{`RANDOM}};
  predictor_114 = _RAND_115[1:0];
  _RAND_116 = {1{`RANDOM}};
  predictor_115 = _RAND_116[1:0];
  _RAND_117 = {1{`RANDOM}};
  predictor_116 = _RAND_117[1:0];
  _RAND_118 = {1{`RANDOM}};
  predictor_117 = _RAND_118[1:0];
  _RAND_119 = {1{`RANDOM}};
  predictor_118 = _RAND_119[1:0];
  _RAND_120 = {1{`RANDOM}};
  predictor_119 = _RAND_120[1:0];
  _RAND_121 = {1{`RANDOM}};
  predictor_120 = _RAND_121[1:0];
  _RAND_122 = {1{`RANDOM}};
  predictor_121 = _RAND_122[1:0];
  _RAND_123 = {1{`RANDOM}};
  predictor_122 = _RAND_123[1:0];
  _RAND_124 = {1{`RANDOM}};
  predictor_123 = _RAND_124[1:0];
  _RAND_125 = {1{`RANDOM}};
  predictor_124 = _RAND_125[1:0];
  _RAND_126 = {1{`RANDOM}};
  predictor_125 = _RAND_126[1:0];
  _RAND_127 = {1{`RANDOM}};
  predictor_126 = _RAND_127[1:0];
  _RAND_128 = {1{`RANDOM}};
  predictor_127 = _RAND_128[1:0];
  _RAND_129 = {1{`RANDOM}};
  bpu_inst_packet_o_data_0 = _RAND_129[31:0];
  _RAND_130 = {1{`RANDOM}};
  bpu_inst_packet_o_data_1 = _RAND_130[31:0];
  _RAND_131 = {1{`RANDOM}};
  bpu_inst_packet_o_data_2 = _RAND_131[31:0];
  _RAND_132 = {1{`RANDOM}};
  bpu_inst_packet_o_data_3 = _RAND_132[31:0];
  _RAND_133 = {1{`RANDOM}};
  bpu_inst_packet_o_data_4 = _RAND_133[31:0];
  _RAND_134 = {1{`RANDOM}};
  bpu_inst_packet_o_data_5 = _RAND_134[31:0];
  _RAND_135 = {1{`RANDOM}};
  bpu_inst_packet_o_data_6 = _RAND_135[31:0];
  _RAND_136 = {1{`RANDOM}};
  bpu_inst_packet_o_data_7 = _RAND_136[31:0];
  _RAND_137 = {1{`RANDOM}};
  bpu_inst_packet_o_addr = _RAND_137[31:0];
  _RAND_138 = {1{`RANDOM}};
  bpu_inst_packet_o_gh_backup = _RAND_138[3:0];
  _RAND_139 = {1{`RANDOM}};
  bpu_inst_packet_o_valid_mask_0 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  bpu_inst_packet_o_valid_mask_1 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  bpu_inst_packet_o_valid_mask_2 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  bpu_inst_packet_o_valid_mask_3 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  bpu_inst_packet_o_valid_mask_4 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  bpu_inst_packet_o_valid_mask_5 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  bpu_inst_packet_o_valid_mask_6 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  bpu_inst_packet_o_valid_mask_7 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  bpu_inst_packet_o_predict_mask_0 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  bpu_inst_packet_o_predict_mask_1 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  bpu_inst_packet_o_predict_mask_2 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  bpu_inst_packet_o_predict_mask_3 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  bpu_inst_packet_o_predict_mask_4 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  bpu_inst_packet_o_predict_mask_5 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  bpu_inst_packet_o_predict_mask_6 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  bpu_inst_packet_o_predict_mask_7 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  bpu_inst_packet_o_valid = _RAND_155[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module ICache(
  input          clock,
  input          reset,
  output         io_icache_req_ready,
  input          io_icache_req_valid,
  input  [31:0]  io_icache_req_bits_addr,
  output         io_icache_resp_valid,
  output [31:0]  io_icache_resp_bits_data_0,
  output [31:0]  io_icache_resp_bits_data_1,
  output [31:0]  io_icache_resp_bits_data_2,
  output [31:0]  io_icache_resp_bits_data_3,
  output [31:0]  io_icache_resp_bits_data_4,
  output [31:0]  io_icache_resp_bits_data_5,
  output [31:0]  io_icache_resp_bits_data_6,
  output [31:0]  io_icache_resp_bits_data_7,
  output [31:0]  io_icache_resp_bits_addr,
  input          io_io_read_req_ready,
  output         io_io_read_req_valid,
  output [31:0]  io_io_read_req_bits_addr,
  input  [255:0] io_io_read_resp_bits_data,
  output         io_icache_debug_state,
  output         io_icache_debug_hit_cache,
  output         io_icache_debug_cache_we,
  output [19:0]  io_icache_debug_cache_read_tag,
  output         io_icache_debug_icache_req_valid,
  output [31:0]  io_icache_debug_icache_req_bits_addr
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_24;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
`endif // RANDOMIZE_REG_INIT
  reg [19:0] cache_tag [0:127]; // @[Icache.scala 54:30]
  wire [19:0] cache_tag_cache_read_tag_MPORT_data; // @[Icache.scala 54:30]
  wire [6:0] cache_tag_cache_read_tag_MPORT_addr; // @[Icache.scala 54:30]
  wire [19:0] cache_tag_MPORT_data; // @[Icache.scala 54:30]
  wire [6:0] cache_tag_MPORT_addr; // @[Icache.scala 54:30]
  wire  cache_tag_MPORT_mask; // @[Icache.scala 54:30]
  wire  cache_tag_MPORT_en; // @[Icache.scala 54:30]
  reg  cache_tag_cache_read_tag_MPORT_en_pipe_0;
  reg [6:0] cache_tag_cache_read_tag_MPORT_addr_pipe_0;
  reg [31:0] cache_data_0 [0:127]; // @[Icache.scala 55:53]
  wire [31:0] cache_data_0_MPORT_9_data; // @[Icache.scala 55:53]
  wire [6:0] cache_data_0_MPORT_9_addr; // @[Icache.scala 55:53]
  wire [31:0] cache_data_0_MPORT_1_data; // @[Icache.scala 55:53]
  wire [6:0] cache_data_0_MPORT_1_addr; // @[Icache.scala 55:53]
  wire  cache_data_0_MPORT_1_mask; // @[Icache.scala 55:53]
  wire  cache_data_0_MPORT_1_en; // @[Icache.scala 55:53]
  reg  cache_data_0_MPORT_9_en_pipe_0;
  reg [6:0] cache_data_0_MPORT_9_addr_pipe_0;
  reg [31:0] cache_data_1 [0:127]; // @[Icache.scala 55:53]
  wire [31:0] cache_data_1_MPORT_10_data; // @[Icache.scala 55:53]
  wire [6:0] cache_data_1_MPORT_10_addr; // @[Icache.scala 55:53]
  wire [31:0] cache_data_1_MPORT_2_data; // @[Icache.scala 55:53]
  wire [6:0] cache_data_1_MPORT_2_addr; // @[Icache.scala 55:53]
  wire  cache_data_1_MPORT_2_mask; // @[Icache.scala 55:53]
  wire  cache_data_1_MPORT_2_en; // @[Icache.scala 55:53]
  reg  cache_data_1_MPORT_10_en_pipe_0;
  reg [6:0] cache_data_1_MPORT_10_addr_pipe_0;
  reg [31:0] cache_data_2 [0:127]; // @[Icache.scala 55:53]
  wire [31:0] cache_data_2_MPORT_11_data; // @[Icache.scala 55:53]
  wire [6:0] cache_data_2_MPORT_11_addr; // @[Icache.scala 55:53]
  wire [31:0] cache_data_2_MPORT_3_data; // @[Icache.scala 55:53]
  wire [6:0] cache_data_2_MPORT_3_addr; // @[Icache.scala 55:53]
  wire  cache_data_2_MPORT_3_mask; // @[Icache.scala 55:53]
  wire  cache_data_2_MPORT_3_en; // @[Icache.scala 55:53]
  reg  cache_data_2_MPORT_11_en_pipe_0;
  reg [6:0] cache_data_2_MPORT_11_addr_pipe_0;
  reg [31:0] cache_data_3 [0:127]; // @[Icache.scala 55:53]
  wire [31:0] cache_data_3_MPORT_12_data; // @[Icache.scala 55:53]
  wire [6:0] cache_data_3_MPORT_12_addr; // @[Icache.scala 55:53]
  wire [31:0] cache_data_3_MPORT_4_data; // @[Icache.scala 55:53]
  wire [6:0] cache_data_3_MPORT_4_addr; // @[Icache.scala 55:53]
  wire  cache_data_3_MPORT_4_mask; // @[Icache.scala 55:53]
  wire  cache_data_3_MPORT_4_en; // @[Icache.scala 55:53]
  reg  cache_data_3_MPORT_12_en_pipe_0;
  reg [6:0] cache_data_3_MPORT_12_addr_pipe_0;
  reg [31:0] cache_data_4 [0:127]; // @[Icache.scala 55:53]
  wire [31:0] cache_data_4_MPORT_13_data; // @[Icache.scala 55:53]
  wire [6:0] cache_data_4_MPORT_13_addr; // @[Icache.scala 55:53]
  wire [31:0] cache_data_4_MPORT_5_data; // @[Icache.scala 55:53]
  wire [6:0] cache_data_4_MPORT_5_addr; // @[Icache.scala 55:53]
  wire  cache_data_4_MPORT_5_mask; // @[Icache.scala 55:53]
  wire  cache_data_4_MPORT_5_en; // @[Icache.scala 55:53]
  reg  cache_data_4_MPORT_13_en_pipe_0;
  reg [6:0] cache_data_4_MPORT_13_addr_pipe_0;
  reg [31:0] cache_data_5 [0:127]; // @[Icache.scala 55:53]
  wire [31:0] cache_data_5_MPORT_14_data; // @[Icache.scala 55:53]
  wire [6:0] cache_data_5_MPORT_14_addr; // @[Icache.scala 55:53]
  wire [31:0] cache_data_5_MPORT_6_data; // @[Icache.scala 55:53]
  wire [6:0] cache_data_5_MPORT_6_addr; // @[Icache.scala 55:53]
  wire  cache_data_5_MPORT_6_mask; // @[Icache.scala 55:53]
  wire  cache_data_5_MPORT_6_en; // @[Icache.scala 55:53]
  reg  cache_data_5_MPORT_14_en_pipe_0;
  reg [6:0] cache_data_5_MPORT_14_addr_pipe_0;
  reg [31:0] cache_data_6 [0:127]; // @[Icache.scala 55:53]
  wire [31:0] cache_data_6_MPORT_15_data; // @[Icache.scala 55:53]
  wire [6:0] cache_data_6_MPORT_15_addr; // @[Icache.scala 55:53]
  wire [31:0] cache_data_6_MPORT_7_data; // @[Icache.scala 55:53]
  wire [6:0] cache_data_6_MPORT_7_addr; // @[Icache.scala 55:53]
  wire  cache_data_6_MPORT_7_mask; // @[Icache.scala 55:53]
  wire  cache_data_6_MPORT_7_en; // @[Icache.scala 55:53]
  reg  cache_data_6_MPORT_15_en_pipe_0;
  reg [6:0] cache_data_6_MPORT_15_addr_pipe_0;
  reg [31:0] cache_data_7 [0:127]; // @[Icache.scala 55:53]
  wire [31:0] cache_data_7_MPORT_16_data; // @[Icache.scala 55:53]
  wire [6:0] cache_data_7_MPORT_16_addr; // @[Icache.scala 55:53]
  wire [31:0] cache_data_7_MPORT_8_data; // @[Icache.scala 55:53]
  wire [6:0] cache_data_7_MPORT_8_addr; // @[Icache.scala 55:53]
  wire  cache_data_7_MPORT_8_mask; // @[Icache.scala 55:53]
  wire  cache_data_7_MPORT_8_en; // @[Icache.scala 55:53]
  reg  cache_data_7_MPORT_16_en_pipe_0;
  reg [6:0] cache_data_7_MPORT_16_addr_pipe_0;
  reg  state; // @[Icache.scala 52:22]
  reg  cache_valid_0; // @[Icache.scala 53:28]
  reg  cache_valid_1; // @[Icache.scala 53:28]
  reg  cache_valid_2; // @[Icache.scala 53:28]
  reg  cache_valid_3; // @[Icache.scala 53:28]
  reg  cache_valid_4; // @[Icache.scala 53:28]
  reg  cache_valid_5; // @[Icache.scala 53:28]
  reg  cache_valid_6; // @[Icache.scala 53:28]
  reg  cache_valid_7; // @[Icache.scala 53:28]
  reg  cache_valid_8; // @[Icache.scala 53:28]
  reg  cache_valid_9; // @[Icache.scala 53:28]
  reg  cache_valid_10; // @[Icache.scala 53:28]
  reg  cache_valid_11; // @[Icache.scala 53:28]
  reg  cache_valid_12; // @[Icache.scala 53:28]
  reg  cache_valid_13; // @[Icache.scala 53:28]
  reg  cache_valid_14; // @[Icache.scala 53:28]
  reg  cache_valid_15; // @[Icache.scala 53:28]
  reg  cache_valid_16; // @[Icache.scala 53:28]
  reg  cache_valid_17; // @[Icache.scala 53:28]
  reg  cache_valid_18; // @[Icache.scala 53:28]
  reg  cache_valid_19; // @[Icache.scala 53:28]
  reg  cache_valid_20; // @[Icache.scala 53:28]
  reg  cache_valid_21; // @[Icache.scala 53:28]
  reg  cache_valid_22; // @[Icache.scala 53:28]
  reg  cache_valid_23; // @[Icache.scala 53:28]
  reg  cache_valid_24; // @[Icache.scala 53:28]
  reg  cache_valid_25; // @[Icache.scala 53:28]
  reg  cache_valid_26; // @[Icache.scala 53:28]
  reg  cache_valid_27; // @[Icache.scala 53:28]
  reg  cache_valid_28; // @[Icache.scala 53:28]
  reg  cache_valid_29; // @[Icache.scala 53:28]
  reg  cache_valid_30; // @[Icache.scala 53:28]
  reg  cache_valid_31; // @[Icache.scala 53:28]
  reg  cache_valid_32; // @[Icache.scala 53:28]
  reg  cache_valid_33; // @[Icache.scala 53:28]
  reg  cache_valid_34; // @[Icache.scala 53:28]
  reg  cache_valid_35; // @[Icache.scala 53:28]
  reg  cache_valid_36; // @[Icache.scala 53:28]
  reg  cache_valid_37; // @[Icache.scala 53:28]
  reg  cache_valid_38; // @[Icache.scala 53:28]
  reg  cache_valid_39; // @[Icache.scala 53:28]
  reg  cache_valid_40; // @[Icache.scala 53:28]
  reg  cache_valid_41; // @[Icache.scala 53:28]
  reg  cache_valid_42; // @[Icache.scala 53:28]
  reg  cache_valid_43; // @[Icache.scala 53:28]
  reg  cache_valid_44; // @[Icache.scala 53:28]
  reg  cache_valid_45; // @[Icache.scala 53:28]
  reg  cache_valid_46; // @[Icache.scala 53:28]
  reg  cache_valid_47; // @[Icache.scala 53:28]
  reg  cache_valid_48; // @[Icache.scala 53:28]
  reg  cache_valid_49; // @[Icache.scala 53:28]
  reg  cache_valid_50; // @[Icache.scala 53:28]
  reg  cache_valid_51; // @[Icache.scala 53:28]
  reg  cache_valid_52; // @[Icache.scala 53:28]
  reg  cache_valid_53; // @[Icache.scala 53:28]
  reg  cache_valid_54; // @[Icache.scala 53:28]
  reg  cache_valid_55; // @[Icache.scala 53:28]
  reg  cache_valid_56; // @[Icache.scala 53:28]
  reg  cache_valid_57; // @[Icache.scala 53:28]
  reg  cache_valid_58; // @[Icache.scala 53:28]
  reg  cache_valid_59; // @[Icache.scala 53:28]
  reg  cache_valid_60; // @[Icache.scala 53:28]
  reg  cache_valid_61; // @[Icache.scala 53:28]
  reg  cache_valid_62; // @[Icache.scala 53:28]
  reg  cache_valid_63; // @[Icache.scala 53:28]
  reg  cache_valid_64; // @[Icache.scala 53:28]
  reg  cache_valid_65; // @[Icache.scala 53:28]
  reg  cache_valid_66; // @[Icache.scala 53:28]
  reg  cache_valid_67; // @[Icache.scala 53:28]
  reg  cache_valid_68; // @[Icache.scala 53:28]
  reg  cache_valid_69; // @[Icache.scala 53:28]
  reg  cache_valid_70; // @[Icache.scala 53:28]
  reg  cache_valid_71; // @[Icache.scala 53:28]
  reg  cache_valid_72; // @[Icache.scala 53:28]
  reg  cache_valid_73; // @[Icache.scala 53:28]
  reg  cache_valid_74; // @[Icache.scala 53:28]
  reg  cache_valid_75; // @[Icache.scala 53:28]
  reg  cache_valid_76; // @[Icache.scala 53:28]
  reg  cache_valid_77; // @[Icache.scala 53:28]
  reg  cache_valid_78; // @[Icache.scala 53:28]
  reg  cache_valid_79; // @[Icache.scala 53:28]
  reg  cache_valid_80; // @[Icache.scala 53:28]
  reg  cache_valid_81; // @[Icache.scala 53:28]
  reg  cache_valid_82; // @[Icache.scala 53:28]
  reg  cache_valid_83; // @[Icache.scala 53:28]
  reg  cache_valid_84; // @[Icache.scala 53:28]
  reg  cache_valid_85; // @[Icache.scala 53:28]
  reg  cache_valid_86; // @[Icache.scala 53:28]
  reg  cache_valid_87; // @[Icache.scala 53:28]
  reg  cache_valid_88; // @[Icache.scala 53:28]
  reg  cache_valid_89; // @[Icache.scala 53:28]
  reg  cache_valid_90; // @[Icache.scala 53:28]
  reg  cache_valid_91; // @[Icache.scala 53:28]
  reg  cache_valid_92; // @[Icache.scala 53:28]
  reg  cache_valid_93; // @[Icache.scala 53:28]
  reg  cache_valid_94; // @[Icache.scala 53:28]
  reg  cache_valid_95; // @[Icache.scala 53:28]
  reg  cache_valid_96; // @[Icache.scala 53:28]
  reg  cache_valid_97; // @[Icache.scala 53:28]
  reg  cache_valid_98; // @[Icache.scala 53:28]
  reg  cache_valid_99; // @[Icache.scala 53:28]
  reg  cache_valid_100; // @[Icache.scala 53:28]
  reg  cache_valid_101; // @[Icache.scala 53:28]
  reg  cache_valid_102; // @[Icache.scala 53:28]
  reg  cache_valid_103; // @[Icache.scala 53:28]
  reg  cache_valid_104; // @[Icache.scala 53:28]
  reg  cache_valid_105; // @[Icache.scala 53:28]
  reg  cache_valid_106; // @[Icache.scala 53:28]
  reg  cache_valid_107; // @[Icache.scala 53:28]
  reg  cache_valid_108; // @[Icache.scala 53:28]
  reg  cache_valid_109; // @[Icache.scala 53:28]
  reg  cache_valid_110; // @[Icache.scala 53:28]
  reg  cache_valid_111; // @[Icache.scala 53:28]
  reg  cache_valid_112; // @[Icache.scala 53:28]
  reg  cache_valid_113; // @[Icache.scala 53:28]
  reg  cache_valid_114; // @[Icache.scala 53:28]
  reg  cache_valid_115; // @[Icache.scala 53:28]
  reg  cache_valid_116; // @[Icache.scala 53:28]
  reg  cache_valid_117; // @[Icache.scala 53:28]
  reg  cache_valid_118; // @[Icache.scala 53:28]
  reg  cache_valid_119; // @[Icache.scala 53:28]
  reg  cache_valid_120; // @[Icache.scala 53:28]
  reg  cache_valid_121; // @[Icache.scala 53:28]
  reg  cache_valid_122; // @[Icache.scala 53:28]
  reg  cache_valid_123; // @[Icache.scala 53:28]
  reg  cache_valid_124; // @[Icache.scala 53:28]
  reg  cache_valid_125; // @[Icache.scala 53:28]
  reg  cache_valid_126; // @[Icache.scala 53:28]
  reg  cache_valid_127; // @[Icache.scala 53:28]
  wire [31:0] io_read_data_0 = io_io_read_resp_bits_data[31:0]; // @[Icache.scala 56:56]
  wire [31:0] io_read_data_1 = io_io_read_resp_bits_data[63:32]; // @[Icache.scala 56:56]
  wire [31:0] io_read_data_2 = io_io_read_resp_bits_data[95:64]; // @[Icache.scala 56:56]
  wire [31:0] io_read_data_3 = io_io_read_resp_bits_data[127:96]; // @[Icache.scala 56:56]
  wire [31:0] io_read_data_4 = io_io_read_resp_bits_data[159:128]; // @[Icache.scala 56:56]
  wire [31:0] io_read_data_5 = io_io_read_resp_bits_data[191:160]; // @[Icache.scala 56:56]
  wire [31:0] io_read_data_6 = io_io_read_resp_bits_data[223:192]; // @[Icache.scala 56:56]
  wire [31:0] io_read_data_7 = io_io_read_resp_bits_data[255:224]; // @[Icache.scala 56:56]
  wire  _T = ~state; // @[Conditional.scala 37:30]
  wire  _GEN_185 = state & io_io_read_req_ready; // @[Conditional.scala 39:67 Icache.scala 72:12]
  wire  cache_we = _T ? 1'h0 : _GEN_185; // @[Conditional.scala 40:58 Icache.scala 72:12]
  wire [19:0] cache_read_tag = cache_tag_cache_read_tag_MPORT_data; // @[Icache.scala 122:19 Icache.scala 128:22]
  wire  _GEN_1 = 7'h1 == io_icache_req_bits_addr[11:5] ? cache_valid_1 : cache_valid_0; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_2 = 7'h2 == io_icache_req_bits_addr[11:5] ? cache_valid_2 : _GEN_1; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_3 = 7'h3 == io_icache_req_bits_addr[11:5] ? cache_valid_3 : _GEN_2; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_4 = 7'h4 == io_icache_req_bits_addr[11:5] ? cache_valid_4 : _GEN_3; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_5 = 7'h5 == io_icache_req_bits_addr[11:5] ? cache_valid_5 : _GEN_4; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_6 = 7'h6 == io_icache_req_bits_addr[11:5] ? cache_valid_6 : _GEN_5; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_7 = 7'h7 == io_icache_req_bits_addr[11:5] ? cache_valid_7 : _GEN_6; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_8 = 7'h8 == io_icache_req_bits_addr[11:5] ? cache_valid_8 : _GEN_7; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_9 = 7'h9 == io_icache_req_bits_addr[11:5] ? cache_valid_9 : _GEN_8; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_10 = 7'ha == io_icache_req_bits_addr[11:5] ? cache_valid_10 : _GEN_9; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_11 = 7'hb == io_icache_req_bits_addr[11:5] ? cache_valid_11 : _GEN_10; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_12 = 7'hc == io_icache_req_bits_addr[11:5] ? cache_valid_12 : _GEN_11; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_13 = 7'hd == io_icache_req_bits_addr[11:5] ? cache_valid_13 : _GEN_12; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_14 = 7'he == io_icache_req_bits_addr[11:5] ? cache_valid_14 : _GEN_13; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_15 = 7'hf == io_icache_req_bits_addr[11:5] ? cache_valid_15 : _GEN_14; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_16 = 7'h10 == io_icache_req_bits_addr[11:5] ? cache_valid_16 : _GEN_15; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_17 = 7'h11 == io_icache_req_bits_addr[11:5] ? cache_valid_17 : _GEN_16; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_18 = 7'h12 == io_icache_req_bits_addr[11:5] ? cache_valid_18 : _GEN_17; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_19 = 7'h13 == io_icache_req_bits_addr[11:5] ? cache_valid_19 : _GEN_18; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_20 = 7'h14 == io_icache_req_bits_addr[11:5] ? cache_valid_20 : _GEN_19; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_21 = 7'h15 == io_icache_req_bits_addr[11:5] ? cache_valid_21 : _GEN_20; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_22 = 7'h16 == io_icache_req_bits_addr[11:5] ? cache_valid_22 : _GEN_21; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_23 = 7'h17 == io_icache_req_bits_addr[11:5] ? cache_valid_23 : _GEN_22; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_24 = 7'h18 == io_icache_req_bits_addr[11:5] ? cache_valid_24 : _GEN_23; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_25 = 7'h19 == io_icache_req_bits_addr[11:5] ? cache_valid_25 : _GEN_24; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_26 = 7'h1a == io_icache_req_bits_addr[11:5] ? cache_valid_26 : _GEN_25; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_27 = 7'h1b == io_icache_req_bits_addr[11:5] ? cache_valid_27 : _GEN_26; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_28 = 7'h1c == io_icache_req_bits_addr[11:5] ? cache_valid_28 : _GEN_27; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_29 = 7'h1d == io_icache_req_bits_addr[11:5] ? cache_valid_29 : _GEN_28; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_30 = 7'h1e == io_icache_req_bits_addr[11:5] ? cache_valid_30 : _GEN_29; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_31 = 7'h1f == io_icache_req_bits_addr[11:5] ? cache_valid_31 : _GEN_30; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_32 = 7'h20 == io_icache_req_bits_addr[11:5] ? cache_valid_32 : _GEN_31; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_33 = 7'h21 == io_icache_req_bits_addr[11:5] ? cache_valid_33 : _GEN_32; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_34 = 7'h22 == io_icache_req_bits_addr[11:5] ? cache_valid_34 : _GEN_33; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_35 = 7'h23 == io_icache_req_bits_addr[11:5] ? cache_valid_35 : _GEN_34; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_36 = 7'h24 == io_icache_req_bits_addr[11:5] ? cache_valid_36 : _GEN_35; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_37 = 7'h25 == io_icache_req_bits_addr[11:5] ? cache_valid_37 : _GEN_36; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_38 = 7'h26 == io_icache_req_bits_addr[11:5] ? cache_valid_38 : _GEN_37; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_39 = 7'h27 == io_icache_req_bits_addr[11:5] ? cache_valid_39 : _GEN_38; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_40 = 7'h28 == io_icache_req_bits_addr[11:5] ? cache_valid_40 : _GEN_39; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_41 = 7'h29 == io_icache_req_bits_addr[11:5] ? cache_valid_41 : _GEN_40; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_42 = 7'h2a == io_icache_req_bits_addr[11:5] ? cache_valid_42 : _GEN_41; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_43 = 7'h2b == io_icache_req_bits_addr[11:5] ? cache_valid_43 : _GEN_42; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_44 = 7'h2c == io_icache_req_bits_addr[11:5] ? cache_valid_44 : _GEN_43; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_45 = 7'h2d == io_icache_req_bits_addr[11:5] ? cache_valid_45 : _GEN_44; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_46 = 7'h2e == io_icache_req_bits_addr[11:5] ? cache_valid_46 : _GEN_45; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_47 = 7'h2f == io_icache_req_bits_addr[11:5] ? cache_valid_47 : _GEN_46; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_48 = 7'h30 == io_icache_req_bits_addr[11:5] ? cache_valid_48 : _GEN_47; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_49 = 7'h31 == io_icache_req_bits_addr[11:5] ? cache_valid_49 : _GEN_48; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_50 = 7'h32 == io_icache_req_bits_addr[11:5] ? cache_valid_50 : _GEN_49; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_51 = 7'h33 == io_icache_req_bits_addr[11:5] ? cache_valid_51 : _GEN_50; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_52 = 7'h34 == io_icache_req_bits_addr[11:5] ? cache_valid_52 : _GEN_51; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_53 = 7'h35 == io_icache_req_bits_addr[11:5] ? cache_valid_53 : _GEN_52; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_54 = 7'h36 == io_icache_req_bits_addr[11:5] ? cache_valid_54 : _GEN_53; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_55 = 7'h37 == io_icache_req_bits_addr[11:5] ? cache_valid_55 : _GEN_54; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_56 = 7'h38 == io_icache_req_bits_addr[11:5] ? cache_valid_56 : _GEN_55; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_57 = 7'h39 == io_icache_req_bits_addr[11:5] ? cache_valid_57 : _GEN_56; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_58 = 7'h3a == io_icache_req_bits_addr[11:5] ? cache_valid_58 : _GEN_57; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_59 = 7'h3b == io_icache_req_bits_addr[11:5] ? cache_valid_59 : _GEN_58; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_60 = 7'h3c == io_icache_req_bits_addr[11:5] ? cache_valid_60 : _GEN_59; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_61 = 7'h3d == io_icache_req_bits_addr[11:5] ? cache_valid_61 : _GEN_60; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_62 = 7'h3e == io_icache_req_bits_addr[11:5] ? cache_valid_62 : _GEN_61; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_63 = 7'h3f == io_icache_req_bits_addr[11:5] ? cache_valid_63 : _GEN_62; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_64 = 7'h40 == io_icache_req_bits_addr[11:5] ? cache_valid_64 : _GEN_63; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_65 = 7'h41 == io_icache_req_bits_addr[11:5] ? cache_valid_65 : _GEN_64; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_66 = 7'h42 == io_icache_req_bits_addr[11:5] ? cache_valid_66 : _GEN_65; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_67 = 7'h43 == io_icache_req_bits_addr[11:5] ? cache_valid_67 : _GEN_66; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_68 = 7'h44 == io_icache_req_bits_addr[11:5] ? cache_valid_68 : _GEN_67; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_69 = 7'h45 == io_icache_req_bits_addr[11:5] ? cache_valid_69 : _GEN_68; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_70 = 7'h46 == io_icache_req_bits_addr[11:5] ? cache_valid_70 : _GEN_69; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_71 = 7'h47 == io_icache_req_bits_addr[11:5] ? cache_valid_71 : _GEN_70; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_72 = 7'h48 == io_icache_req_bits_addr[11:5] ? cache_valid_72 : _GEN_71; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_73 = 7'h49 == io_icache_req_bits_addr[11:5] ? cache_valid_73 : _GEN_72; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_74 = 7'h4a == io_icache_req_bits_addr[11:5] ? cache_valid_74 : _GEN_73; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_75 = 7'h4b == io_icache_req_bits_addr[11:5] ? cache_valid_75 : _GEN_74; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_76 = 7'h4c == io_icache_req_bits_addr[11:5] ? cache_valid_76 : _GEN_75; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_77 = 7'h4d == io_icache_req_bits_addr[11:5] ? cache_valid_77 : _GEN_76; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_78 = 7'h4e == io_icache_req_bits_addr[11:5] ? cache_valid_78 : _GEN_77; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_79 = 7'h4f == io_icache_req_bits_addr[11:5] ? cache_valid_79 : _GEN_78; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_80 = 7'h50 == io_icache_req_bits_addr[11:5] ? cache_valid_80 : _GEN_79; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_81 = 7'h51 == io_icache_req_bits_addr[11:5] ? cache_valid_81 : _GEN_80; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_82 = 7'h52 == io_icache_req_bits_addr[11:5] ? cache_valid_82 : _GEN_81; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_83 = 7'h53 == io_icache_req_bits_addr[11:5] ? cache_valid_83 : _GEN_82; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_84 = 7'h54 == io_icache_req_bits_addr[11:5] ? cache_valid_84 : _GEN_83; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_85 = 7'h55 == io_icache_req_bits_addr[11:5] ? cache_valid_85 : _GEN_84; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_86 = 7'h56 == io_icache_req_bits_addr[11:5] ? cache_valid_86 : _GEN_85; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_87 = 7'h57 == io_icache_req_bits_addr[11:5] ? cache_valid_87 : _GEN_86; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_88 = 7'h58 == io_icache_req_bits_addr[11:5] ? cache_valid_88 : _GEN_87; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_89 = 7'h59 == io_icache_req_bits_addr[11:5] ? cache_valid_89 : _GEN_88; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_90 = 7'h5a == io_icache_req_bits_addr[11:5] ? cache_valid_90 : _GEN_89; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_91 = 7'h5b == io_icache_req_bits_addr[11:5] ? cache_valid_91 : _GEN_90; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_92 = 7'h5c == io_icache_req_bits_addr[11:5] ? cache_valid_92 : _GEN_91; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_93 = 7'h5d == io_icache_req_bits_addr[11:5] ? cache_valid_93 : _GEN_92; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_94 = 7'h5e == io_icache_req_bits_addr[11:5] ? cache_valid_94 : _GEN_93; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_95 = 7'h5f == io_icache_req_bits_addr[11:5] ? cache_valid_95 : _GEN_94; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_96 = 7'h60 == io_icache_req_bits_addr[11:5] ? cache_valid_96 : _GEN_95; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_97 = 7'h61 == io_icache_req_bits_addr[11:5] ? cache_valid_97 : _GEN_96; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_98 = 7'h62 == io_icache_req_bits_addr[11:5] ? cache_valid_98 : _GEN_97; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_99 = 7'h63 == io_icache_req_bits_addr[11:5] ? cache_valid_99 : _GEN_98; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_100 = 7'h64 == io_icache_req_bits_addr[11:5] ? cache_valid_100 : _GEN_99; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_101 = 7'h65 == io_icache_req_bits_addr[11:5] ? cache_valid_101 : _GEN_100; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_102 = 7'h66 == io_icache_req_bits_addr[11:5] ? cache_valid_102 : _GEN_101; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_103 = 7'h67 == io_icache_req_bits_addr[11:5] ? cache_valid_103 : _GEN_102; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_104 = 7'h68 == io_icache_req_bits_addr[11:5] ? cache_valid_104 : _GEN_103; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_105 = 7'h69 == io_icache_req_bits_addr[11:5] ? cache_valid_105 : _GEN_104; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_106 = 7'h6a == io_icache_req_bits_addr[11:5] ? cache_valid_106 : _GEN_105; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_107 = 7'h6b == io_icache_req_bits_addr[11:5] ? cache_valid_107 : _GEN_106; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_108 = 7'h6c == io_icache_req_bits_addr[11:5] ? cache_valid_108 : _GEN_107; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_109 = 7'h6d == io_icache_req_bits_addr[11:5] ? cache_valid_109 : _GEN_108; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_110 = 7'h6e == io_icache_req_bits_addr[11:5] ? cache_valid_110 : _GEN_109; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_111 = 7'h6f == io_icache_req_bits_addr[11:5] ? cache_valid_111 : _GEN_110; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_112 = 7'h70 == io_icache_req_bits_addr[11:5] ? cache_valid_112 : _GEN_111; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_113 = 7'h71 == io_icache_req_bits_addr[11:5] ? cache_valid_113 : _GEN_112; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_114 = 7'h72 == io_icache_req_bits_addr[11:5] ? cache_valid_114 : _GEN_113; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_115 = 7'h73 == io_icache_req_bits_addr[11:5] ? cache_valid_115 : _GEN_114; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_116 = 7'h74 == io_icache_req_bits_addr[11:5] ? cache_valid_116 : _GEN_115; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_117 = 7'h75 == io_icache_req_bits_addr[11:5] ? cache_valid_117 : _GEN_116; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_118 = 7'h76 == io_icache_req_bits_addr[11:5] ? cache_valid_118 : _GEN_117; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_119 = 7'h77 == io_icache_req_bits_addr[11:5] ? cache_valid_119 : _GEN_118; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_120 = 7'h78 == io_icache_req_bits_addr[11:5] ? cache_valid_120 : _GEN_119; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_121 = 7'h79 == io_icache_req_bits_addr[11:5] ? cache_valid_121 : _GEN_120; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_122 = 7'h7a == io_icache_req_bits_addr[11:5] ? cache_valid_122 : _GEN_121; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_123 = 7'h7b == io_icache_req_bits_addr[11:5] ? cache_valid_123 : _GEN_122; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_124 = 7'h7c == io_icache_req_bits_addr[11:5] ? cache_valid_124 : _GEN_123; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_125 = 7'h7d == io_icache_req_bits_addr[11:5] ? cache_valid_125 : _GEN_124; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_126 = 7'h7e == io_icache_req_bits_addr[11:5] ? cache_valid_126 : _GEN_125; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  _GEN_127 = 7'h7f == io_icache_req_bits_addr[11:5] ? cache_valid_127 : _GEN_126; // @[Icache.scala 79:78 Icache.scala 79:78]
  wire  hit_cache = cache_read_tag == io_icache_req_bits_addr[31:12] & _GEN_127; // @[Icache.scala 79:78]
  wire  _GEN_129 = io_icache_req_valid | state; // @[Icache.scala 82:32 Icache.scala 84:14 Icache.scala 52:22]
  wire  _GEN_130 = hit_cache ? 1'h0 : 1'h1; // @[Icache.scala 107:28 Icache.scala 108:29 Icache.scala 115:29]
  wire [31:0] cache_read_data_0 = cache_data_0_MPORT_9_data; // @[Icache.scala 129:33 Icache.scala 129:33]
  wire [31:0] cache_read_data_1 = cache_data_1_MPORT_10_data; // @[Icache.scala 129:33 Icache.scala 129:33]
  wire [31:0] cache_read_data_2 = cache_data_2_MPORT_11_data; // @[Icache.scala 129:33 Icache.scala 129:33]
  wire [31:0] cache_read_data_3 = cache_data_3_MPORT_12_data; // @[Icache.scala 129:33 Icache.scala 129:33]
  wire [31:0] cache_read_data_4 = cache_data_4_MPORT_13_data; // @[Icache.scala 129:33 Icache.scala 129:33]
  wire [31:0] cache_read_data_5 = cache_data_5_MPORT_14_data; // @[Icache.scala 129:33 Icache.scala 129:33]
  wire [31:0] cache_read_data_6 = cache_data_6_MPORT_15_data; // @[Icache.scala 129:33 Icache.scala 129:33]
  wire [31:0] cache_read_data_7 = cache_data_7_MPORT_16_data; // @[Icache.scala 129:33 Icache.scala 129:33]
  wire  _GEN_140 = hit_cache ? 1'h0 : state; // @[Icache.scala 107:28 Icache.scala 113:14 Icache.scala 52:22]
  wire  _GEN_141 = ~io_icache_req_valid ? 1'h0 : _GEN_130; // @[Icache.scala 101:39 Icache.scala 102:29]
  wire  _GEN_150 = ~io_icache_req_valid ? 1'h0 : hit_cache; // @[Icache.scala 101:39 Icache.scala 104:29]
  wire  _GEN_151 = ~io_icache_req_valid ? 1'h0 : _GEN_140; // @[Icache.scala 101:39 Icache.scala 106:14]
  wire  _GEN_152 = io_io_read_req_ready ? 1'h0 : _GEN_141; // @[Icache.scala 90:33 Icache.scala 91:29]
  wire  _GEN_153 = io_io_read_req_ready ? io_icache_req_valid : _GEN_150; // @[Icache.scala 90:33 Icache.scala 92:29]
  wire  _GEN_162 = io_io_read_req_ready | _GEN_150; // @[Icache.scala 90:33 Icache.scala 94:28]
  wire [19:0] _GEN_164 = io_io_read_req_ready ? io_icache_req_bits_addr[31:12] : 20'h0; // @[Icache.scala 90:33 Icache.scala 97:24 Icache.scala 77:19]
  wire [31:0] _GEN_165 = io_io_read_req_ready ? io_read_data_0 : 32'h0; // @[Icache.scala 90:33 Icache.scala 98:25 Icache.scala 78:20]
  wire [31:0] _GEN_166 = io_io_read_req_ready ? io_read_data_1 : 32'h0; // @[Icache.scala 90:33 Icache.scala 98:25 Icache.scala 78:20]
  wire [31:0] _GEN_167 = io_io_read_req_ready ? io_read_data_2 : 32'h0; // @[Icache.scala 90:33 Icache.scala 98:25 Icache.scala 78:20]
  wire [31:0] _GEN_168 = io_io_read_req_ready ? io_read_data_3 : 32'h0; // @[Icache.scala 90:33 Icache.scala 98:25 Icache.scala 78:20]
  wire [31:0] _GEN_169 = io_io_read_req_ready ? io_read_data_4 : 32'h0; // @[Icache.scala 90:33 Icache.scala 98:25 Icache.scala 78:20]
  wire [31:0] _GEN_170 = io_io_read_req_ready ? io_read_data_5 : 32'h0; // @[Icache.scala 90:33 Icache.scala 98:25 Icache.scala 78:20]
  wire [31:0] _GEN_171 = io_io_read_req_ready ? io_read_data_6 : 32'h0; // @[Icache.scala 90:33 Icache.scala 98:25 Icache.scala 78:20]
  wire [31:0] _GEN_172 = io_io_read_req_ready ? io_read_data_7 : 32'h0; // @[Icache.scala 90:33 Icache.scala 98:25 Icache.scala 78:20]
  wire  _GEN_174 = state & _GEN_152; // @[Conditional.scala 39:67 Icache.scala 67:23]
  wire  _GEN_175 = state & _GEN_153; // @[Conditional.scala 39:67 Icache.scala 70:23]
  wire  _GEN_184 = state & _GEN_162; // @[Conditional.scala 39:67 Icache.scala 68:22]
  wire [19:0] _GEN_186 = state ? _GEN_164 : 20'h0; // @[Conditional.scala 39:67 Icache.scala 77:19]
  wire [31:0] _GEN_187 = state ? _GEN_165 : 32'h0; // @[Conditional.scala 39:67 Icache.scala 78:20]
  wire [31:0] _GEN_188 = state ? _GEN_166 : 32'h0; // @[Conditional.scala 39:67 Icache.scala 78:20]
  wire [31:0] _GEN_189 = state ? _GEN_167 : 32'h0; // @[Conditional.scala 39:67 Icache.scala 78:20]
  wire [31:0] _GEN_190 = state ? _GEN_168 : 32'h0; // @[Conditional.scala 39:67 Icache.scala 78:20]
  wire [31:0] _GEN_191 = state ? _GEN_169 : 32'h0; // @[Conditional.scala 39:67 Icache.scala 78:20]
  wire [31:0] _GEN_192 = state ? _GEN_170 : 32'h0; // @[Conditional.scala 39:67 Icache.scala 78:20]
  wire [31:0] _GEN_193 = state ? _GEN_171 : 32'h0; // @[Conditional.scala 39:67 Icache.scala 78:20]
  wire [31:0] _GEN_194 = state ? _GEN_172 : 32'h0; // @[Conditional.scala 39:67 Icache.scala 78:20]
  wire  _GEN_300 = 7'h0 == io_icache_req_bits_addr[11:5] | cache_valid_0; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_301 = 7'h1 == io_icache_req_bits_addr[11:5] | cache_valid_1; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_302 = 7'h2 == io_icache_req_bits_addr[11:5] | cache_valid_2; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_303 = 7'h3 == io_icache_req_bits_addr[11:5] | cache_valid_3; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_304 = 7'h4 == io_icache_req_bits_addr[11:5] | cache_valid_4; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_305 = 7'h5 == io_icache_req_bits_addr[11:5] | cache_valid_5; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_306 = 7'h6 == io_icache_req_bits_addr[11:5] | cache_valid_6; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_307 = 7'h7 == io_icache_req_bits_addr[11:5] | cache_valid_7; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_308 = 7'h8 == io_icache_req_bits_addr[11:5] | cache_valid_8; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_309 = 7'h9 == io_icache_req_bits_addr[11:5] | cache_valid_9; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_310 = 7'ha == io_icache_req_bits_addr[11:5] | cache_valid_10; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_311 = 7'hb == io_icache_req_bits_addr[11:5] | cache_valid_11; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_312 = 7'hc == io_icache_req_bits_addr[11:5] | cache_valid_12; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_313 = 7'hd == io_icache_req_bits_addr[11:5] | cache_valid_13; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_314 = 7'he == io_icache_req_bits_addr[11:5] | cache_valid_14; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_315 = 7'hf == io_icache_req_bits_addr[11:5] | cache_valid_15; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_316 = 7'h10 == io_icache_req_bits_addr[11:5] | cache_valid_16; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_317 = 7'h11 == io_icache_req_bits_addr[11:5] | cache_valid_17; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_318 = 7'h12 == io_icache_req_bits_addr[11:5] | cache_valid_18; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_319 = 7'h13 == io_icache_req_bits_addr[11:5] | cache_valid_19; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_320 = 7'h14 == io_icache_req_bits_addr[11:5] | cache_valid_20; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_321 = 7'h15 == io_icache_req_bits_addr[11:5] | cache_valid_21; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_322 = 7'h16 == io_icache_req_bits_addr[11:5] | cache_valid_22; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_323 = 7'h17 == io_icache_req_bits_addr[11:5] | cache_valid_23; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_324 = 7'h18 == io_icache_req_bits_addr[11:5] | cache_valid_24; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_325 = 7'h19 == io_icache_req_bits_addr[11:5] | cache_valid_25; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_326 = 7'h1a == io_icache_req_bits_addr[11:5] | cache_valid_26; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_327 = 7'h1b == io_icache_req_bits_addr[11:5] | cache_valid_27; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_328 = 7'h1c == io_icache_req_bits_addr[11:5] | cache_valid_28; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_329 = 7'h1d == io_icache_req_bits_addr[11:5] | cache_valid_29; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_330 = 7'h1e == io_icache_req_bits_addr[11:5] | cache_valid_30; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_331 = 7'h1f == io_icache_req_bits_addr[11:5] | cache_valid_31; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_332 = 7'h20 == io_icache_req_bits_addr[11:5] | cache_valid_32; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_333 = 7'h21 == io_icache_req_bits_addr[11:5] | cache_valid_33; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_334 = 7'h22 == io_icache_req_bits_addr[11:5] | cache_valid_34; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_335 = 7'h23 == io_icache_req_bits_addr[11:5] | cache_valid_35; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_336 = 7'h24 == io_icache_req_bits_addr[11:5] | cache_valid_36; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_337 = 7'h25 == io_icache_req_bits_addr[11:5] | cache_valid_37; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_338 = 7'h26 == io_icache_req_bits_addr[11:5] | cache_valid_38; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_339 = 7'h27 == io_icache_req_bits_addr[11:5] | cache_valid_39; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_340 = 7'h28 == io_icache_req_bits_addr[11:5] | cache_valid_40; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_341 = 7'h29 == io_icache_req_bits_addr[11:5] | cache_valid_41; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_342 = 7'h2a == io_icache_req_bits_addr[11:5] | cache_valid_42; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_343 = 7'h2b == io_icache_req_bits_addr[11:5] | cache_valid_43; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_344 = 7'h2c == io_icache_req_bits_addr[11:5] | cache_valid_44; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_345 = 7'h2d == io_icache_req_bits_addr[11:5] | cache_valid_45; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_346 = 7'h2e == io_icache_req_bits_addr[11:5] | cache_valid_46; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_347 = 7'h2f == io_icache_req_bits_addr[11:5] | cache_valid_47; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_348 = 7'h30 == io_icache_req_bits_addr[11:5] | cache_valid_48; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_349 = 7'h31 == io_icache_req_bits_addr[11:5] | cache_valid_49; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_350 = 7'h32 == io_icache_req_bits_addr[11:5] | cache_valid_50; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_351 = 7'h33 == io_icache_req_bits_addr[11:5] | cache_valid_51; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_352 = 7'h34 == io_icache_req_bits_addr[11:5] | cache_valid_52; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_353 = 7'h35 == io_icache_req_bits_addr[11:5] | cache_valid_53; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_354 = 7'h36 == io_icache_req_bits_addr[11:5] | cache_valid_54; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_355 = 7'h37 == io_icache_req_bits_addr[11:5] | cache_valid_55; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_356 = 7'h38 == io_icache_req_bits_addr[11:5] | cache_valid_56; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_357 = 7'h39 == io_icache_req_bits_addr[11:5] | cache_valid_57; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_358 = 7'h3a == io_icache_req_bits_addr[11:5] | cache_valid_58; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_359 = 7'h3b == io_icache_req_bits_addr[11:5] | cache_valid_59; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_360 = 7'h3c == io_icache_req_bits_addr[11:5] | cache_valid_60; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_361 = 7'h3d == io_icache_req_bits_addr[11:5] | cache_valid_61; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_362 = 7'h3e == io_icache_req_bits_addr[11:5] | cache_valid_62; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_363 = 7'h3f == io_icache_req_bits_addr[11:5] | cache_valid_63; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_364 = 7'h40 == io_icache_req_bits_addr[11:5] | cache_valid_64; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_365 = 7'h41 == io_icache_req_bits_addr[11:5] | cache_valid_65; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_366 = 7'h42 == io_icache_req_bits_addr[11:5] | cache_valid_66; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_367 = 7'h43 == io_icache_req_bits_addr[11:5] | cache_valid_67; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_368 = 7'h44 == io_icache_req_bits_addr[11:5] | cache_valid_68; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_369 = 7'h45 == io_icache_req_bits_addr[11:5] | cache_valid_69; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_370 = 7'h46 == io_icache_req_bits_addr[11:5] | cache_valid_70; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_371 = 7'h47 == io_icache_req_bits_addr[11:5] | cache_valid_71; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_372 = 7'h48 == io_icache_req_bits_addr[11:5] | cache_valid_72; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_373 = 7'h49 == io_icache_req_bits_addr[11:5] | cache_valid_73; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_374 = 7'h4a == io_icache_req_bits_addr[11:5] | cache_valid_74; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_375 = 7'h4b == io_icache_req_bits_addr[11:5] | cache_valid_75; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_376 = 7'h4c == io_icache_req_bits_addr[11:5] | cache_valid_76; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_377 = 7'h4d == io_icache_req_bits_addr[11:5] | cache_valid_77; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_378 = 7'h4e == io_icache_req_bits_addr[11:5] | cache_valid_78; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_379 = 7'h4f == io_icache_req_bits_addr[11:5] | cache_valid_79; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_380 = 7'h50 == io_icache_req_bits_addr[11:5] | cache_valid_80; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_381 = 7'h51 == io_icache_req_bits_addr[11:5] | cache_valid_81; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_382 = 7'h52 == io_icache_req_bits_addr[11:5] | cache_valid_82; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_383 = 7'h53 == io_icache_req_bits_addr[11:5] | cache_valid_83; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_384 = 7'h54 == io_icache_req_bits_addr[11:5] | cache_valid_84; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_385 = 7'h55 == io_icache_req_bits_addr[11:5] | cache_valid_85; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_386 = 7'h56 == io_icache_req_bits_addr[11:5] | cache_valid_86; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_387 = 7'h57 == io_icache_req_bits_addr[11:5] | cache_valid_87; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_388 = 7'h58 == io_icache_req_bits_addr[11:5] | cache_valid_88; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_389 = 7'h59 == io_icache_req_bits_addr[11:5] | cache_valid_89; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_390 = 7'h5a == io_icache_req_bits_addr[11:5] | cache_valid_90; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_391 = 7'h5b == io_icache_req_bits_addr[11:5] | cache_valid_91; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_392 = 7'h5c == io_icache_req_bits_addr[11:5] | cache_valid_92; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_393 = 7'h5d == io_icache_req_bits_addr[11:5] | cache_valid_93; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_394 = 7'h5e == io_icache_req_bits_addr[11:5] | cache_valid_94; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_395 = 7'h5f == io_icache_req_bits_addr[11:5] | cache_valid_95; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_396 = 7'h60 == io_icache_req_bits_addr[11:5] | cache_valid_96; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_397 = 7'h61 == io_icache_req_bits_addr[11:5] | cache_valid_97; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_398 = 7'h62 == io_icache_req_bits_addr[11:5] | cache_valid_98; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_399 = 7'h63 == io_icache_req_bits_addr[11:5] | cache_valid_99; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_400 = 7'h64 == io_icache_req_bits_addr[11:5] | cache_valid_100; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_401 = 7'h65 == io_icache_req_bits_addr[11:5] | cache_valid_101; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_402 = 7'h66 == io_icache_req_bits_addr[11:5] | cache_valid_102; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_403 = 7'h67 == io_icache_req_bits_addr[11:5] | cache_valid_103; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_404 = 7'h68 == io_icache_req_bits_addr[11:5] | cache_valid_104; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_405 = 7'h69 == io_icache_req_bits_addr[11:5] | cache_valid_105; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_406 = 7'h6a == io_icache_req_bits_addr[11:5] | cache_valid_106; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_407 = 7'h6b == io_icache_req_bits_addr[11:5] | cache_valid_107; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_408 = 7'h6c == io_icache_req_bits_addr[11:5] | cache_valid_108; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_409 = 7'h6d == io_icache_req_bits_addr[11:5] | cache_valid_109; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_410 = 7'h6e == io_icache_req_bits_addr[11:5] | cache_valid_110; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_411 = 7'h6f == io_icache_req_bits_addr[11:5] | cache_valid_111; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_412 = 7'h70 == io_icache_req_bits_addr[11:5] | cache_valid_112; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_413 = 7'h71 == io_icache_req_bits_addr[11:5] | cache_valid_113; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_414 = 7'h72 == io_icache_req_bits_addr[11:5] | cache_valid_114; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_415 = 7'h73 == io_icache_req_bits_addr[11:5] | cache_valid_115; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_416 = 7'h74 == io_icache_req_bits_addr[11:5] | cache_valid_116; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_417 = 7'h75 == io_icache_req_bits_addr[11:5] | cache_valid_117; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_418 = 7'h76 == io_icache_req_bits_addr[11:5] | cache_valid_118; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_419 = 7'h77 == io_icache_req_bits_addr[11:5] | cache_valid_119; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_420 = 7'h78 == io_icache_req_bits_addr[11:5] | cache_valid_120; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_421 = 7'h79 == io_icache_req_bits_addr[11:5] | cache_valid_121; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_422 = 7'h7a == io_icache_req_bits_addr[11:5] | cache_valid_122; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_423 = 7'h7b == io_icache_req_bits_addr[11:5] | cache_valid_123; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_424 = 7'h7c == io_icache_req_bits_addr[11:5] | cache_valid_124; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_425 = 7'h7d == io_icache_req_bits_addr[11:5] | cache_valid_125; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_426 = 7'h7e == io_icache_req_bits_addr[11:5] | cache_valid_126; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire  _GEN_427 = 7'h7f == io_icache_req_bits_addr[11:5] | cache_valid_127; // @[Icache.scala 136:103 Icache.scala 136:103 Icache.scala 53:28]
  wire [26:0] io_io_read_req_bits_addr_hi = io_icache_req_bits_addr[31:5]; // @[Icache.scala 139:58]
  assign cache_tag_cache_read_tag_MPORT_addr = cache_tag_cache_read_tag_MPORT_addr_pipe_0;
  assign cache_tag_cache_read_tag_MPORT_data = cache_tag[cache_tag_cache_read_tag_MPORT_addr]; // @[Icache.scala 54:30]
  assign cache_tag_MPORT_data = _T ? 20'h0 : _GEN_186;
  assign cache_tag_MPORT_addr = io_icache_req_bits_addr[11:5];
  assign cache_tag_MPORT_mask = 1'h1;
  assign cache_tag_MPORT_en = _T ? 1'h0 : _GEN_185;
  assign cache_data_0_MPORT_9_addr = cache_data_0_MPORT_9_addr_pipe_0;
  assign cache_data_0_MPORT_9_data = cache_data_0[cache_data_0_MPORT_9_addr]; // @[Icache.scala 55:53]
  assign cache_data_0_MPORT_1_data = _T ? 32'h0 : _GEN_187;
  assign cache_data_0_MPORT_1_addr = io_icache_req_bits_addr[11:5];
  assign cache_data_0_MPORT_1_mask = 1'h1;
  assign cache_data_0_MPORT_1_en = _T ? 1'h0 : _GEN_185;
  assign cache_data_1_MPORT_10_addr = cache_data_1_MPORT_10_addr_pipe_0;
  assign cache_data_1_MPORT_10_data = cache_data_1[cache_data_1_MPORT_10_addr]; // @[Icache.scala 55:53]
  assign cache_data_1_MPORT_2_data = _T ? 32'h0 : _GEN_188;
  assign cache_data_1_MPORT_2_addr = io_icache_req_bits_addr[11:5];
  assign cache_data_1_MPORT_2_mask = 1'h1;
  assign cache_data_1_MPORT_2_en = _T ? 1'h0 : _GEN_185;
  assign cache_data_2_MPORT_11_addr = cache_data_2_MPORT_11_addr_pipe_0;
  assign cache_data_2_MPORT_11_data = cache_data_2[cache_data_2_MPORT_11_addr]; // @[Icache.scala 55:53]
  assign cache_data_2_MPORT_3_data = _T ? 32'h0 : _GEN_189;
  assign cache_data_2_MPORT_3_addr = io_icache_req_bits_addr[11:5];
  assign cache_data_2_MPORT_3_mask = 1'h1;
  assign cache_data_2_MPORT_3_en = _T ? 1'h0 : _GEN_185;
  assign cache_data_3_MPORT_12_addr = cache_data_3_MPORT_12_addr_pipe_0;
  assign cache_data_3_MPORT_12_data = cache_data_3[cache_data_3_MPORT_12_addr]; // @[Icache.scala 55:53]
  assign cache_data_3_MPORT_4_data = _T ? 32'h0 : _GEN_190;
  assign cache_data_3_MPORT_4_addr = io_icache_req_bits_addr[11:5];
  assign cache_data_3_MPORT_4_mask = 1'h1;
  assign cache_data_3_MPORT_4_en = _T ? 1'h0 : _GEN_185;
  assign cache_data_4_MPORT_13_addr = cache_data_4_MPORT_13_addr_pipe_0;
  assign cache_data_4_MPORT_13_data = cache_data_4[cache_data_4_MPORT_13_addr]; // @[Icache.scala 55:53]
  assign cache_data_4_MPORT_5_data = _T ? 32'h0 : _GEN_191;
  assign cache_data_4_MPORT_5_addr = io_icache_req_bits_addr[11:5];
  assign cache_data_4_MPORT_5_mask = 1'h1;
  assign cache_data_4_MPORT_5_en = _T ? 1'h0 : _GEN_185;
  assign cache_data_5_MPORT_14_addr = cache_data_5_MPORT_14_addr_pipe_0;
  assign cache_data_5_MPORT_14_data = cache_data_5[cache_data_5_MPORT_14_addr]; // @[Icache.scala 55:53]
  assign cache_data_5_MPORT_6_data = _T ? 32'h0 : _GEN_192;
  assign cache_data_5_MPORT_6_addr = io_icache_req_bits_addr[11:5];
  assign cache_data_5_MPORT_6_mask = 1'h1;
  assign cache_data_5_MPORT_6_en = _T ? 1'h0 : _GEN_185;
  assign cache_data_6_MPORT_15_addr = cache_data_6_MPORT_15_addr_pipe_0;
  assign cache_data_6_MPORT_15_data = cache_data_6[cache_data_6_MPORT_15_addr]; // @[Icache.scala 55:53]
  assign cache_data_6_MPORT_7_data = _T ? 32'h0 : _GEN_193;
  assign cache_data_6_MPORT_7_addr = io_icache_req_bits_addr[11:5];
  assign cache_data_6_MPORT_7_mask = 1'h1;
  assign cache_data_6_MPORT_7_en = _T ? 1'h0 : _GEN_185;
  assign cache_data_7_MPORT_16_addr = cache_data_7_MPORT_16_addr_pipe_0;
  assign cache_data_7_MPORT_16_data = cache_data_7[cache_data_7_MPORT_16_addr]; // @[Icache.scala 55:53]
  assign cache_data_7_MPORT_8_data = _T ? 32'h0 : _GEN_194;
  assign cache_data_7_MPORT_8_addr = io_icache_req_bits_addr[11:5];
  assign cache_data_7_MPORT_8_mask = 1'h1;
  assign cache_data_7_MPORT_8_en = _T ? 1'h0 : _GEN_185;
  assign io_icache_req_ready = _T ? 1'h0 : _GEN_184; // @[Conditional.scala 40:58 Icache.scala 68:22]
  assign io_icache_resp_valid = _T ? 1'h0 : _GEN_175; // @[Conditional.scala 40:58 Icache.scala 70:23]
  assign io_icache_resp_bits_data_0 = io_io_read_req_ready ? io_read_data_0 : cache_read_data_0; // @[Icache.scala 90:33 Icache.scala 93:33]
  assign io_icache_resp_bits_data_1 = io_io_read_req_ready ? io_read_data_1 : cache_read_data_1; // @[Icache.scala 90:33 Icache.scala 93:33]
  assign io_icache_resp_bits_data_2 = io_io_read_req_ready ? io_read_data_2 : cache_read_data_2; // @[Icache.scala 90:33 Icache.scala 93:33]
  assign io_icache_resp_bits_data_3 = io_io_read_req_ready ? io_read_data_3 : cache_read_data_3; // @[Icache.scala 90:33 Icache.scala 93:33]
  assign io_icache_resp_bits_data_4 = io_io_read_req_ready ? io_read_data_4 : cache_read_data_4; // @[Icache.scala 90:33 Icache.scala 93:33]
  assign io_icache_resp_bits_data_5 = io_io_read_req_ready ? io_read_data_5 : cache_read_data_5; // @[Icache.scala 90:33 Icache.scala 93:33]
  assign io_icache_resp_bits_data_6 = io_io_read_req_ready ? io_read_data_6 : cache_read_data_6; // @[Icache.scala 90:33 Icache.scala 93:33]
  assign io_icache_resp_bits_data_7 = io_io_read_req_ready ? io_read_data_7 : cache_read_data_7; // @[Icache.scala 90:33 Icache.scala 93:33]
  assign io_icache_resp_bits_addr = io_icache_req_bits_addr; // @[Icache.scala 141:27]
  assign io_io_read_req_valid = _T ? io_icache_req_valid : _GEN_174; // @[Conditional.scala 40:58]
  assign io_io_read_req_bits_addr = {io_io_read_req_bits_addr_hi,5'h0}; // @[Cat.scala 30:58]
  assign io_icache_debug_state = state; // @[Icache.scala 147:24]
  assign io_icache_debug_hit_cache = cache_read_tag == io_icache_req_bits_addr[31:12] & _GEN_127; // @[Icache.scala 79:78]
  assign io_icache_debug_cache_we = _T ? 1'h0 : _GEN_185; // @[Conditional.scala 40:58 Icache.scala 72:12]
  assign io_icache_debug_cache_read_tag = cache_tag_cache_read_tag_MPORT_data; // @[Icache.scala 122:19 Icache.scala 128:22]
  assign io_icache_debug_icache_req_valid = io_icache_req_valid; // @[Icache.scala 145:35]
  assign io_icache_debug_icache_req_bits_addr = io_icache_req_bits_addr; // @[Icache.scala 146:39]
  always @(posedge clock) begin
    if(cache_tag_MPORT_en & cache_tag_MPORT_mask) begin
      cache_tag[cache_tag_MPORT_addr] <= cache_tag_MPORT_data; // @[Icache.scala 54:30]
    end
    if (cache_we) begin
      cache_tag_cache_read_tag_MPORT_en_pipe_0 <= 1'h0;
    end else begin
      cache_tag_cache_read_tag_MPORT_en_pipe_0 <= 1'h1;
    end
    if (cache_we ? 1'h0 : 1'h1) begin
      cache_tag_cache_read_tag_MPORT_addr_pipe_0 <= io_icache_req_bits_addr[11:5];
    end
    if(cache_data_0_MPORT_1_en & cache_data_0_MPORT_1_mask) begin
      cache_data_0[cache_data_0_MPORT_1_addr] <= cache_data_0_MPORT_1_data; // @[Icache.scala 55:53]
    end
    if (cache_we) begin
      cache_data_0_MPORT_9_en_pipe_0 <= 1'h0;
    end else begin
      cache_data_0_MPORT_9_en_pipe_0 <= 1'h1;
    end
    if (cache_we ? 1'h0 : 1'h1) begin
      cache_data_0_MPORT_9_addr_pipe_0 <= io_icache_req_bits_addr[11:5];
    end
    if(cache_data_1_MPORT_2_en & cache_data_1_MPORT_2_mask) begin
      cache_data_1[cache_data_1_MPORT_2_addr] <= cache_data_1_MPORT_2_data; // @[Icache.scala 55:53]
    end
    if (cache_we) begin
      cache_data_1_MPORT_10_en_pipe_0 <= 1'h0;
    end else begin
      cache_data_1_MPORT_10_en_pipe_0 <= 1'h1;
    end
    if (cache_we ? 1'h0 : 1'h1) begin
      cache_data_1_MPORT_10_addr_pipe_0 <= io_icache_req_bits_addr[11:5];
    end
    if(cache_data_2_MPORT_3_en & cache_data_2_MPORT_3_mask) begin
      cache_data_2[cache_data_2_MPORT_3_addr] <= cache_data_2_MPORT_3_data; // @[Icache.scala 55:53]
    end
    if (cache_we) begin
      cache_data_2_MPORT_11_en_pipe_0 <= 1'h0;
    end else begin
      cache_data_2_MPORT_11_en_pipe_0 <= 1'h1;
    end
    if (cache_we ? 1'h0 : 1'h1) begin
      cache_data_2_MPORT_11_addr_pipe_0 <= io_icache_req_bits_addr[11:5];
    end
    if(cache_data_3_MPORT_4_en & cache_data_3_MPORT_4_mask) begin
      cache_data_3[cache_data_3_MPORT_4_addr] <= cache_data_3_MPORT_4_data; // @[Icache.scala 55:53]
    end
    if (cache_we) begin
      cache_data_3_MPORT_12_en_pipe_0 <= 1'h0;
    end else begin
      cache_data_3_MPORT_12_en_pipe_0 <= 1'h1;
    end
    if (cache_we ? 1'h0 : 1'h1) begin
      cache_data_3_MPORT_12_addr_pipe_0 <= io_icache_req_bits_addr[11:5];
    end
    if(cache_data_4_MPORT_5_en & cache_data_4_MPORT_5_mask) begin
      cache_data_4[cache_data_4_MPORT_5_addr] <= cache_data_4_MPORT_5_data; // @[Icache.scala 55:53]
    end
    if (cache_we) begin
      cache_data_4_MPORT_13_en_pipe_0 <= 1'h0;
    end else begin
      cache_data_4_MPORT_13_en_pipe_0 <= 1'h1;
    end
    if (cache_we ? 1'h0 : 1'h1) begin
      cache_data_4_MPORT_13_addr_pipe_0 <= io_icache_req_bits_addr[11:5];
    end
    if(cache_data_5_MPORT_6_en & cache_data_5_MPORT_6_mask) begin
      cache_data_5[cache_data_5_MPORT_6_addr] <= cache_data_5_MPORT_6_data; // @[Icache.scala 55:53]
    end
    if (cache_we) begin
      cache_data_5_MPORT_14_en_pipe_0 <= 1'h0;
    end else begin
      cache_data_5_MPORT_14_en_pipe_0 <= 1'h1;
    end
    if (cache_we ? 1'h0 : 1'h1) begin
      cache_data_5_MPORT_14_addr_pipe_0 <= io_icache_req_bits_addr[11:5];
    end
    if(cache_data_6_MPORT_7_en & cache_data_6_MPORT_7_mask) begin
      cache_data_6[cache_data_6_MPORT_7_addr] <= cache_data_6_MPORT_7_data; // @[Icache.scala 55:53]
    end
    if (cache_we) begin
      cache_data_6_MPORT_15_en_pipe_0 <= 1'h0;
    end else begin
      cache_data_6_MPORT_15_en_pipe_0 <= 1'h1;
    end
    if (cache_we ? 1'h0 : 1'h1) begin
      cache_data_6_MPORT_15_addr_pipe_0 <= io_icache_req_bits_addr[11:5];
    end
    if(cache_data_7_MPORT_8_en & cache_data_7_MPORT_8_mask) begin
      cache_data_7[cache_data_7_MPORT_8_addr] <= cache_data_7_MPORT_8_data; // @[Icache.scala 55:53]
    end
    if (cache_we) begin
      cache_data_7_MPORT_16_en_pipe_0 <= 1'h0;
    end else begin
      cache_data_7_MPORT_16_en_pipe_0 <= 1'h1;
    end
    if (cache_we ? 1'h0 : 1'h1) begin
      cache_data_7_MPORT_16_addr_pipe_0 <= io_icache_req_bits_addr[11:5];
    end
    if (reset) begin // @[Icache.scala 52:22]
      state <= 1'h0; // @[Icache.scala 52:22]
    end else if (_T) begin // @[Conditional.scala 40:58]
      state <= _GEN_129;
    end else if (state) begin // @[Conditional.scala 39:67]
      if (io_io_read_req_ready) begin // @[Icache.scala 90:33]
        state <= 1'h0; // @[Icache.scala 100:14]
      end else begin
        state <= _GEN_151;
      end
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_0 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_0 <= _GEN_300;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_1 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_1 <= _GEN_301;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_2 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_2 <= _GEN_302;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_3 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_3 <= _GEN_303;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_4 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_4 <= _GEN_304;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_5 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_5 <= _GEN_305;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_6 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_6 <= _GEN_306;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_7 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_7 <= _GEN_307;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_8 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_8 <= _GEN_308;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_9 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_9 <= _GEN_309;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_10 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_10 <= _GEN_310;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_11 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_11 <= _GEN_311;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_12 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_12 <= _GEN_312;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_13 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_13 <= _GEN_313;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_14 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_14 <= _GEN_314;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_15 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_15 <= _GEN_315;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_16 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_16 <= _GEN_316;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_17 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_17 <= _GEN_317;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_18 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_18 <= _GEN_318;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_19 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_19 <= _GEN_319;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_20 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_20 <= _GEN_320;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_21 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_21 <= _GEN_321;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_22 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_22 <= _GEN_322;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_23 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_23 <= _GEN_323;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_24 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_24 <= _GEN_324;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_25 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_25 <= _GEN_325;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_26 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_26 <= _GEN_326;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_27 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_27 <= _GEN_327;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_28 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_28 <= _GEN_328;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_29 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_29 <= _GEN_329;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_30 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_30 <= _GEN_330;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_31 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_31 <= _GEN_331;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_32 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_32 <= _GEN_332;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_33 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_33 <= _GEN_333;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_34 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_34 <= _GEN_334;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_35 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_35 <= _GEN_335;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_36 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_36 <= _GEN_336;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_37 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_37 <= _GEN_337;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_38 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_38 <= _GEN_338;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_39 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_39 <= _GEN_339;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_40 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_40 <= _GEN_340;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_41 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_41 <= _GEN_341;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_42 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_42 <= _GEN_342;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_43 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_43 <= _GEN_343;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_44 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_44 <= _GEN_344;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_45 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_45 <= _GEN_345;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_46 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_46 <= _GEN_346;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_47 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_47 <= _GEN_347;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_48 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_48 <= _GEN_348;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_49 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_49 <= _GEN_349;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_50 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_50 <= _GEN_350;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_51 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_51 <= _GEN_351;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_52 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_52 <= _GEN_352;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_53 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_53 <= _GEN_353;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_54 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_54 <= _GEN_354;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_55 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_55 <= _GEN_355;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_56 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_56 <= _GEN_356;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_57 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_57 <= _GEN_357;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_58 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_58 <= _GEN_358;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_59 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_59 <= _GEN_359;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_60 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_60 <= _GEN_360;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_61 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_61 <= _GEN_361;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_62 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_62 <= _GEN_362;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_63 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_63 <= _GEN_363;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_64 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_64 <= _GEN_364;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_65 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_65 <= _GEN_365;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_66 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_66 <= _GEN_366;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_67 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_67 <= _GEN_367;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_68 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_68 <= _GEN_368;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_69 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_69 <= _GEN_369;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_70 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_70 <= _GEN_370;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_71 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_71 <= _GEN_371;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_72 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_72 <= _GEN_372;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_73 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_73 <= _GEN_373;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_74 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_74 <= _GEN_374;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_75 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_75 <= _GEN_375;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_76 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_76 <= _GEN_376;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_77 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_77 <= _GEN_377;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_78 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_78 <= _GEN_378;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_79 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_79 <= _GEN_379;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_80 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_80 <= _GEN_380;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_81 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_81 <= _GEN_381;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_82 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_82 <= _GEN_382;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_83 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_83 <= _GEN_383;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_84 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_84 <= _GEN_384;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_85 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_85 <= _GEN_385;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_86 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_86 <= _GEN_386;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_87 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_87 <= _GEN_387;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_88 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_88 <= _GEN_388;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_89 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_89 <= _GEN_389;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_90 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_90 <= _GEN_390;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_91 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_91 <= _GEN_391;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_92 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_92 <= _GEN_392;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_93 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_93 <= _GEN_393;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_94 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_94 <= _GEN_394;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_95 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_95 <= _GEN_395;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_96 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_96 <= _GEN_396;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_97 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_97 <= _GEN_397;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_98 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_98 <= _GEN_398;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_99 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_99 <= _GEN_399;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_100 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_100 <= _GEN_400;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_101 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_101 <= _GEN_401;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_102 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_102 <= _GEN_402;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_103 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_103 <= _GEN_403;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_104 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_104 <= _GEN_404;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_105 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_105 <= _GEN_405;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_106 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_106 <= _GEN_406;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_107 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_107 <= _GEN_407;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_108 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_108 <= _GEN_408;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_109 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_109 <= _GEN_409;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_110 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_110 <= _GEN_410;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_111 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_111 <= _GEN_411;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_112 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_112 <= _GEN_412;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_113 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_113 <= _GEN_413;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_114 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_114 <= _GEN_414;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_115 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_115 <= _GEN_415;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_116 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_116 <= _GEN_416;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_117 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_117 <= _GEN_417;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_118 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_118 <= _GEN_418;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_119 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_119 <= _GEN_419;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_120 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_120 <= _GEN_420;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_121 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_121 <= _GEN_421;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_122 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_122 <= _GEN_422;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_123 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_123 <= _GEN_423;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_124 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_124 <= _GEN_424;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_125 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_125 <= _GEN_425;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_126 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_126 <= _GEN_426;
    end
    if (reset) begin // @[Icache.scala 53:28]
      cache_valid_127 <= 1'h0; // @[Icache.scala 53:28]
    end else if (cache_we) begin // @[Icache.scala 135:23]
      cache_valid_127 <= _GEN_427;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    cache_tag[initvar] = _RAND_0[19:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    cache_data_0[initvar] = _RAND_3[31:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    cache_data_1[initvar] = _RAND_6[31:0];
  _RAND_9 = {1{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    cache_data_2[initvar] = _RAND_9[31:0];
  _RAND_12 = {1{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    cache_data_3[initvar] = _RAND_12[31:0];
  _RAND_15 = {1{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    cache_data_4[initvar] = _RAND_15[31:0];
  _RAND_18 = {1{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    cache_data_5[initvar] = _RAND_18[31:0];
  _RAND_21 = {1{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    cache_data_6[initvar] = _RAND_21[31:0];
  _RAND_24 = {1{`RANDOM}};
  for (initvar = 0; initvar < 128; initvar = initvar+1)
    cache_data_7[initvar] = _RAND_24[31:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  cache_tag_cache_read_tag_MPORT_en_pipe_0 = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  cache_tag_cache_read_tag_MPORT_addr_pipe_0 = _RAND_2[6:0];
  _RAND_4 = {1{`RANDOM}};
  cache_data_0_MPORT_9_en_pipe_0 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  cache_data_0_MPORT_9_addr_pipe_0 = _RAND_5[6:0];
  _RAND_7 = {1{`RANDOM}};
  cache_data_1_MPORT_10_en_pipe_0 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  cache_data_1_MPORT_10_addr_pipe_0 = _RAND_8[6:0];
  _RAND_10 = {1{`RANDOM}};
  cache_data_2_MPORT_11_en_pipe_0 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  cache_data_2_MPORT_11_addr_pipe_0 = _RAND_11[6:0];
  _RAND_13 = {1{`RANDOM}};
  cache_data_3_MPORT_12_en_pipe_0 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  cache_data_3_MPORT_12_addr_pipe_0 = _RAND_14[6:0];
  _RAND_16 = {1{`RANDOM}};
  cache_data_4_MPORT_13_en_pipe_0 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  cache_data_4_MPORT_13_addr_pipe_0 = _RAND_17[6:0];
  _RAND_19 = {1{`RANDOM}};
  cache_data_5_MPORT_14_en_pipe_0 = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  cache_data_5_MPORT_14_addr_pipe_0 = _RAND_20[6:0];
  _RAND_22 = {1{`RANDOM}};
  cache_data_6_MPORT_15_en_pipe_0 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  cache_data_6_MPORT_15_addr_pipe_0 = _RAND_23[6:0];
  _RAND_25 = {1{`RANDOM}};
  cache_data_7_MPORT_16_en_pipe_0 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  cache_data_7_MPORT_16_addr_pipe_0 = _RAND_26[6:0];
  _RAND_27 = {1{`RANDOM}};
  state = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  cache_valid_0 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  cache_valid_1 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  cache_valid_2 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  cache_valid_3 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  cache_valid_4 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  cache_valid_5 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  cache_valid_6 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  cache_valid_7 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  cache_valid_8 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  cache_valid_9 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  cache_valid_10 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  cache_valid_11 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  cache_valid_12 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  cache_valid_13 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  cache_valid_14 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  cache_valid_15 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  cache_valid_16 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  cache_valid_17 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  cache_valid_18 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  cache_valid_19 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  cache_valid_20 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  cache_valid_21 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  cache_valid_22 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  cache_valid_23 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  cache_valid_24 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  cache_valid_25 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  cache_valid_26 = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  cache_valid_27 = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  cache_valid_28 = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  cache_valid_29 = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  cache_valid_30 = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  cache_valid_31 = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  cache_valid_32 = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  cache_valid_33 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  cache_valid_34 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  cache_valid_35 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  cache_valid_36 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  cache_valid_37 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  cache_valid_38 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  cache_valid_39 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  cache_valid_40 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  cache_valid_41 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  cache_valid_42 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  cache_valid_43 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  cache_valid_44 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  cache_valid_45 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  cache_valid_46 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  cache_valid_47 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  cache_valid_48 = _RAND_76[0:0];
  _RAND_77 = {1{`RANDOM}};
  cache_valid_49 = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  cache_valid_50 = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  cache_valid_51 = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  cache_valid_52 = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  cache_valid_53 = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  cache_valid_54 = _RAND_82[0:0];
  _RAND_83 = {1{`RANDOM}};
  cache_valid_55 = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  cache_valid_56 = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  cache_valid_57 = _RAND_85[0:0];
  _RAND_86 = {1{`RANDOM}};
  cache_valid_58 = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  cache_valid_59 = _RAND_87[0:0];
  _RAND_88 = {1{`RANDOM}};
  cache_valid_60 = _RAND_88[0:0];
  _RAND_89 = {1{`RANDOM}};
  cache_valid_61 = _RAND_89[0:0];
  _RAND_90 = {1{`RANDOM}};
  cache_valid_62 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  cache_valid_63 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  cache_valid_64 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  cache_valid_65 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  cache_valid_66 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  cache_valid_67 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  cache_valid_68 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  cache_valid_69 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  cache_valid_70 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  cache_valid_71 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  cache_valid_72 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  cache_valid_73 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  cache_valid_74 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  cache_valid_75 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  cache_valid_76 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  cache_valid_77 = _RAND_105[0:0];
  _RAND_106 = {1{`RANDOM}};
  cache_valid_78 = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  cache_valid_79 = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  cache_valid_80 = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  cache_valid_81 = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  cache_valid_82 = _RAND_110[0:0];
  _RAND_111 = {1{`RANDOM}};
  cache_valid_83 = _RAND_111[0:0];
  _RAND_112 = {1{`RANDOM}};
  cache_valid_84 = _RAND_112[0:0];
  _RAND_113 = {1{`RANDOM}};
  cache_valid_85 = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  cache_valid_86 = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  cache_valid_87 = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  cache_valid_88 = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  cache_valid_89 = _RAND_117[0:0];
  _RAND_118 = {1{`RANDOM}};
  cache_valid_90 = _RAND_118[0:0];
  _RAND_119 = {1{`RANDOM}};
  cache_valid_91 = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  cache_valid_92 = _RAND_120[0:0];
  _RAND_121 = {1{`RANDOM}};
  cache_valid_93 = _RAND_121[0:0];
  _RAND_122 = {1{`RANDOM}};
  cache_valid_94 = _RAND_122[0:0];
  _RAND_123 = {1{`RANDOM}};
  cache_valid_95 = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  cache_valid_96 = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  cache_valid_97 = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  cache_valid_98 = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  cache_valid_99 = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  cache_valid_100 = _RAND_128[0:0];
  _RAND_129 = {1{`RANDOM}};
  cache_valid_101 = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  cache_valid_102 = _RAND_130[0:0];
  _RAND_131 = {1{`RANDOM}};
  cache_valid_103 = _RAND_131[0:0];
  _RAND_132 = {1{`RANDOM}};
  cache_valid_104 = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  cache_valid_105 = _RAND_133[0:0];
  _RAND_134 = {1{`RANDOM}};
  cache_valid_106 = _RAND_134[0:0];
  _RAND_135 = {1{`RANDOM}};
  cache_valid_107 = _RAND_135[0:0];
  _RAND_136 = {1{`RANDOM}};
  cache_valid_108 = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  cache_valid_109 = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  cache_valid_110 = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  cache_valid_111 = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  cache_valid_112 = _RAND_140[0:0];
  _RAND_141 = {1{`RANDOM}};
  cache_valid_113 = _RAND_141[0:0];
  _RAND_142 = {1{`RANDOM}};
  cache_valid_114 = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  cache_valid_115 = _RAND_143[0:0];
  _RAND_144 = {1{`RANDOM}};
  cache_valid_116 = _RAND_144[0:0];
  _RAND_145 = {1{`RANDOM}};
  cache_valid_117 = _RAND_145[0:0];
  _RAND_146 = {1{`RANDOM}};
  cache_valid_118 = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  cache_valid_119 = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  cache_valid_120 = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  cache_valid_121 = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  cache_valid_122 = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  cache_valid_123 = _RAND_151[0:0];
  _RAND_152 = {1{`RANDOM}};
  cache_valid_124 = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  cache_valid_125 = _RAND_153[0:0];
  _RAND_154 = {1{`RANDOM}};
  cache_valid_126 = _RAND_154[0:0];
  _RAND_155 = {1{`RANDOM}};
  cache_valid_127 = _RAND_155[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module FetchBuffer(
  input         clock,
  input         reset,
  output        io_bpu_inst_packet_i_ready,
  input         io_bpu_inst_packet_i_valid,
  input  [31:0] io_bpu_inst_packet_i_bits_data_0,
  input  [31:0] io_bpu_inst_packet_i_bits_data_1,
  input  [31:0] io_bpu_inst_packet_i_bits_data_2,
  input  [31:0] io_bpu_inst_packet_i_bits_data_3,
  input  [31:0] io_bpu_inst_packet_i_bits_data_4,
  input  [31:0] io_bpu_inst_packet_i_bits_data_5,
  input  [31:0] io_bpu_inst_packet_i_bits_data_6,
  input  [31:0] io_bpu_inst_packet_i_bits_data_7,
  input  [31:0] io_bpu_inst_packet_i_bits_addr,
  input  [3:0]  io_bpu_inst_packet_i_bits_gh_backup,
  input         io_bpu_inst_packet_i_bits_valid_mask_0,
  input         io_bpu_inst_packet_i_bits_valid_mask_1,
  input         io_bpu_inst_packet_i_bits_valid_mask_2,
  input         io_bpu_inst_packet_i_bits_valid_mask_3,
  input         io_bpu_inst_packet_i_bits_valid_mask_4,
  input         io_bpu_inst_packet_i_bits_valid_mask_5,
  input         io_bpu_inst_packet_i_bits_valid_mask_6,
  input         io_bpu_inst_packet_i_bits_valid_mask_7,
  input         io_bpu_inst_packet_i_bits_predict_mask_0,
  input         io_bpu_inst_packet_i_bits_predict_mask_1,
  input         io_bpu_inst_packet_i_bits_predict_mask_2,
  input         io_bpu_inst_packet_i_bits_predict_mask_3,
  input         io_bpu_inst_packet_i_bits_predict_mask_4,
  input         io_bpu_inst_packet_i_bits_predict_mask_5,
  input         io_bpu_inst_packet_i_bits_predict_mask_6,
  input         io_bpu_inst_packet_i_bits_predict_mask_7,
  output        io_inst_bank_valid,
  output [31:0] io_inst_bank_bits_data_0_inst,
  output [31:0] io_inst_bank_bits_data_0_inst_addr,
  output [3:0]  io_inst_bank_bits_data_0_gh_backup,
  output        io_inst_bank_bits_data_0_is_valid,
  output        io_inst_bank_bits_data_0_predict_taken,
  output [31:0] io_inst_bank_bits_data_1_inst,
  output [31:0] io_inst_bank_bits_data_1_inst_addr,
  output [3:0]  io_inst_bank_bits_data_1_gh_backup,
  output        io_inst_bank_bits_data_1_is_valid,
  output        io_inst_bank_bits_data_1_predict_taken,
  input         io_fb_resp_deq_valid_0,
  input         io_fb_resp_deq_valid_1,
  input         io_clear_i
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] fetch_buffer_0_inst; // @[FetchBuffer.scala 50:25]
  reg [31:0] fetch_buffer_0_inst_addr; // @[FetchBuffer.scala 50:25]
  reg [3:0] fetch_buffer_0_gh_backup; // @[FetchBuffer.scala 50:25]
  reg  fetch_buffer_0_predict_taken; // @[FetchBuffer.scala 50:25]
  reg [31:0] fetch_buffer_1_inst; // @[FetchBuffer.scala 50:25]
  reg [31:0] fetch_buffer_1_inst_addr; // @[FetchBuffer.scala 50:25]
  reg [3:0] fetch_buffer_1_gh_backup; // @[FetchBuffer.scala 50:25]
  reg  fetch_buffer_1_predict_taken; // @[FetchBuffer.scala 50:25]
  reg [31:0] fetch_buffer_2_inst; // @[FetchBuffer.scala 50:25]
  reg [31:0] fetch_buffer_2_inst_addr; // @[FetchBuffer.scala 50:25]
  reg [3:0] fetch_buffer_2_gh_backup; // @[FetchBuffer.scala 50:25]
  reg  fetch_buffer_2_predict_taken; // @[FetchBuffer.scala 50:25]
  reg [31:0] fetch_buffer_3_inst; // @[FetchBuffer.scala 50:25]
  reg [31:0] fetch_buffer_3_inst_addr; // @[FetchBuffer.scala 50:25]
  reg [3:0] fetch_buffer_3_gh_backup; // @[FetchBuffer.scala 50:25]
  reg  fetch_buffer_3_predict_taken; // @[FetchBuffer.scala 50:25]
  reg [31:0] fetch_buffer_4_inst; // @[FetchBuffer.scala 50:25]
  reg [31:0] fetch_buffer_4_inst_addr; // @[FetchBuffer.scala 50:25]
  reg [3:0] fetch_buffer_4_gh_backup; // @[FetchBuffer.scala 50:25]
  reg  fetch_buffer_4_predict_taken; // @[FetchBuffer.scala 50:25]
  reg [31:0] fetch_buffer_5_inst; // @[FetchBuffer.scala 50:25]
  reg [31:0] fetch_buffer_5_inst_addr; // @[FetchBuffer.scala 50:25]
  reg [3:0] fetch_buffer_5_gh_backup; // @[FetchBuffer.scala 50:25]
  reg  fetch_buffer_5_predict_taken; // @[FetchBuffer.scala 50:25]
  reg [31:0] fetch_buffer_6_inst; // @[FetchBuffer.scala 50:25]
  reg [31:0] fetch_buffer_6_inst_addr; // @[FetchBuffer.scala 50:25]
  reg [3:0] fetch_buffer_6_gh_backup; // @[FetchBuffer.scala 50:25]
  reg  fetch_buffer_6_predict_taken; // @[FetchBuffer.scala 50:25]
  reg [31:0] fetch_buffer_7_inst; // @[FetchBuffer.scala 50:25]
  reg [31:0] fetch_buffer_7_inst_addr; // @[FetchBuffer.scala 50:25]
  reg [3:0] fetch_buffer_7_gh_backup; // @[FetchBuffer.scala 50:25]
  reg  fetch_buffer_7_predict_taken; // @[FetchBuffer.scala 50:25]
  reg [31:0] fetch_buffer_8_inst; // @[FetchBuffer.scala 50:25]
  reg [31:0] fetch_buffer_8_inst_addr; // @[FetchBuffer.scala 50:25]
  reg [3:0] fetch_buffer_8_gh_backup; // @[FetchBuffer.scala 50:25]
  reg  fetch_buffer_8_predict_taken; // @[FetchBuffer.scala 50:25]
  reg [31:0] fetch_buffer_9_inst; // @[FetchBuffer.scala 50:25]
  reg [31:0] fetch_buffer_9_inst_addr; // @[FetchBuffer.scala 50:25]
  reg [3:0] fetch_buffer_9_gh_backup; // @[FetchBuffer.scala 50:25]
  reg  fetch_buffer_9_predict_taken; // @[FetchBuffer.scala 50:25]
  reg [31:0] fetch_buffer_10_inst; // @[FetchBuffer.scala 50:25]
  reg [31:0] fetch_buffer_10_inst_addr; // @[FetchBuffer.scala 50:25]
  reg [3:0] fetch_buffer_10_gh_backup; // @[FetchBuffer.scala 50:25]
  reg  fetch_buffer_10_predict_taken; // @[FetchBuffer.scala 50:25]
  reg [31:0] fetch_buffer_11_inst; // @[FetchBuffer.scala 50:25]
  reg [31:0] fetch_buffer_11_inst_addr; // @[FetchBuffer.scala 50:25]
  reg [3:0] fetch_buffer_11_gh_backup; // @[FetchBuffer.scala 50:25]
  reg  fetch_buffer_11_predict_taken; // @[FetchBuffer.scala 50:25]
  reg [31:0] fetch_buffer_12_inst; // @[FetchBuffer.scala 50:25]
  reg [31:0] fetch_buffer_12_inst_addr; // @[FetchBuffer.scala 50:25]
  reg [3:0] fetch_buffer_12_gh_backup; // @[FetchBuffer.scala 50:25]
  reg  fetch_buffer_12_predict_taken; // @[FetchBuffer.scala 50:25]
  reg [31:0] fetch_buffer_13_inst; // @[FetchBuffer.scala 50:25]
  reg [31:0] fetch_buffer_13_inst_addr; // @[FetchBuffer.scala 50:25]
  reg [3:0] fetch_buffer_13_gh_backup; // @[FetchBuffer.scala 50:25]
  reg  fetch_buffer_13_predict_taken; // @[FetchBuffer.scala 50:25]
  reg [31:0] fetch_buffer_14_inst; // @[FetchBuffer.scala 50:25]
  reg [31:0] fetch_buffer_14_inst_addr; // @[FetchBuffer.scala 50:25]
  reg [3:0] fetch_buffer_14_gh_backup; // @[FetchBuffer.scala 50:25]
  reg  fetch_buffer_14_predict_taken; // @[FetchBuffer.scala 50:25]
  reg [31:0] fetch_buffer_15_inst; // @[FetchBuffer.scala 50:25]
  reg [31:0] fetch_buffer_15_inst_addr; // @[FetchBuffer.scala 50:25]
  reg [3:0] fetch_buffer_15_gh_backup; // @[FetchBuffer.scala 50:25]
  reg  fetch_buffer_15_predict_taken; // @[FetchBuffer.scala 50:25]
  reg [31:0] fetch_buffer_16_inst; // @[FetchBuffer.scala 50:25]
  reg [31:0] fetch_buffer_16_inst_addr; // @[FetchBuffer.scala 50:25]
  reg [3:0] fetch_buffer_16_gh_backup; // @[FetchBuffer.scala 50:25]
  reg  fetch_buffer_16_predict_taken; // @[FetchBuffer.scala 50:25]
  reg [16:0] deq_idxs_0; // @[FetchBuffer.scala 51:29]
  reg [16:0] tail; // @[FetchBuffer.scala 52:29]
  reg  maybe_full; // @[FetchBuffer.scala 53:29]
  wire  hit_head = deq_idxs_0 == tail; // @[FetchBuffer.scala 55:27]
  wire  is_full = hit_head & maybe_full; // @[FetchBuffer.scala 56:31]
  wire  is_empty = hit_head & ~maybe_full; // @[FetchBuffer.scala 57:31]
  wire [15:0] hi = tail[15:0]; // @[FetchBuffer.scala 42:12]
  wire  lo = tail[16]; // @[FetchBuffer.scala 42:29]
  wire [16:0] _T = {hi,lo}; // @[Cat.scala 30:58]
  wire [16:0] enq_idxs_1 = io_bpu_inst_packet_i_bits_valid_mask_0 ? _T : tail; // @[FetchBuffer.scala 68:18]
  wire [15:0] hi_1 = enq_idxs_1[15:0]; // @[FetchBuffer.scala 42:12]
  wire  lo_1 = enq_idxs_1[16]; // @[FetchBuffer.scala 42:29]
  wire [16:0] _T_2 = {hi_1,lo_1}; // @[Cat.scala 30:58]
  wire [16:0] enq_idxs_2 = io_bpu_inst_packet_i_bits_valid_mask_1 ? _T_2 : enq_idxs_1; // @[FetchBuffer.scala 68:18]
  wire [15:0] hi_2 = enq_idxs_2[15:0]; // @[FetchBuffer.scala 42:12]
  wire  lo_2 = enq_idxs_2[16]; // @[FetchBuffer.scala 42:29]
  wire [16:0] _T_4 = {hi_2,lo_2}; // @[Cat.scala 30:58]
  wire [16:0] enq_idxs_3 = io_bpu_inst_packet_i_bits_valid_mask_2 ? _T_4 : enq_idxs_2; // @[FetchBuffer.scala 68:18]
  wire [15:0] hi_3 = enq_idxs_3[15:0]; // @[FetchBuffer.scala 42:12]
  wire  lo_3 = enq_idxs_3[16]; // @[FetchBuffer.scala 42:29]
  wire [16:0] _T_6 = {hi_3,lo_3}; // @[Cat.scala 30:58]
  wire [16:0] enq_idxs_4 = io_bpu_inst_packet_i_bits_valid_mask_3 ? _T_6 : enq_idxs_3; // @[FetchBuffer.scala 68:18]
  wire [15:0] hi_4 = enq_idxs_4[15:0]; // @[FetchBuffer.scala 42:12]
  wire  lo_4 = enq_idxs_4[16]; // @[FetchBuffer.scala 42:29]
  wire [16:0] _T_8 = {hi_4,lo_4}; // @[Cat.scala 30:58]
  wire [16:0] enq_idxs_5 = io_bpu_inst_packet_i_bits_valid_mask_4 ? _T_8 : enq_idxs_4; // @[FetchBuffer.scala 68:18]
  wire [15:0] hi_5 = enq_idxs_5[15:0]; // @[FetchBuffer.scala 42:12]
  wire  lo_5 = enq_idxs_5[16]; // @[FetchBuffer.scala 42:29]
  wire [16:0] _T_10 = {hi_5,lo_5}; // @[Cat.scala 30:58]
  wire [16:0] enq_idxs_6 = io_bpu_inst_packet_i_bits_valid_mask_5 ? _T_10 : enq_idxs_5; // @[FetchBuffer.scala 68:18]
  wire [15:0] hi_6 = enq_idxs_6[15:0]; // @[FetchBuffer.scala 42:12]
  wire  lo_6 = enq_idxs_6[16]; // @[FetchBuffer.scala 42:29]
  wire [16:0] _T_12 = {hi_6,lo_6}; // @[Cat.scala 30:58]
  wire [16:0] enq_idxs_7 = io_bpu_inst_packet_i_bits_valid_mask_6 ? _T_12 : enq_idxs_6; // @[FetchBuffer.scala 68:18]
  wire  might_hit_head = tail == deq_idxs_0 | enq_idxs_1 == deq_idxs_0 | enq_idxs_2 == deq_idxs_0 | enq_idxs_3 ==
    deq_idxs_0 | enq_idxs_4 == deq_idxs_0 | enq_idxs_5 == deq_idxs_0 | enq_idxs_6 == deq_idxs_0 | enq_idxs_7 ==
    deq_idxs_0; // @[FetchBuffer.scala 61:58]
  wire  _do_enq_T_2 = is_empty | ~(is_full | might_hit_head); // @[FetchBuffer.scala 63:34]
  wire  _do_enq_T_10 = io_bpu_inst_packet_i_bits_valid_mask_0 | io_bpu_inst_packet_i_bits_valid_mask_1 |
    io_bpu_inst_packet_i_bits_valid_mask_2 | io_bpu_inst_packet_i_bits_valid_mask_3 |
    io_bpu_inst_packet_i_bits_valid_mask_4 | io_bpu_inst_packet_i_bits_valid_mask_5 |
    io_bpu_inst_packet_i_bits_valid_mask_6 | io_bpu_inst_packet_i_bits_valid_mask_7; // @[FetchBuffer.scala 63:146]
  wire  do_enq = (is_empty | ~(is_full | might_hit_head)) & io_bpu_inst_packet_i_valid & (
    io_bpu_inst_packet_i_bits_valid_mask_0 | io_bpu_inst_packet_i_bits_valid_mask_1 |
    io_bpu_inst_packet_i_bits_valid_mask_2 | io_bpu_inst_packet_i_bits_valid_mask_3 |
    io_bpu_inst_packet_i_bits_valid_mask_4 | io_bpu_inst_packet_i_bits_valid_mask_5 |
    io_bpu_inst_packet_i_bits_valid_mask_6 | io_bpu_inst_packet_i_bits_valid_mask_7); // @[FetchBuffer.scala 63:97]
  wire [15:0] hi_7 = enq_idxs_7[15:0]; // @[FetchBuffer.scala 42:12]
  wire  lo_7 = enq_idxs_7[16]; // @[FetchBuffer.scala 42:29]
  wire [16:0] _T_14 = {hi_7,lo_7}; // @[Cat.scala 30:58]
  wire [26:0] inst_packet_0_inst_addr_hi_hi = io_bpu_inst_packet_i_bits_addr[31:5]; // @[FetchBuffer.scala 74:67]
  wire [31:0] inst_packet_0_inst_addr = {inst_packet_0_inst_addr_hi_hi,3'h0,2'h0}; // @[Cat.scala 30:58]
  wire [31:0] inst_packet_1_inst_addr = {inst_packet_0_inst_addr_hi_hi,3'h1,2'h0}; // @[Cat.scala 30:58]
  wire [31:0] inst_packet_2_inst_addr = {inst_packet_0_inst_addr_hi_hi,3'h2,2'h0}; // @[Cat.scala 30:58]
  wire [31:0] inst_packet_3_inst_addr = {inst_packet_0_inst_addr_hi_hi,3'h3,2'h0}; // @[Cat.scala 30:58]
  wire [31:0] inst_packet_4_inst_addr = {inst_packet_0_inst_addr_hi_hi,3'h4,2'h0}; // @[Cat.scala 30:58]
  wire [31:0] inst_packet_5_inst_addr = {inst_packet_0_inst_addr_hi_hi,3'h5,2'h0}; // @[Cat.scala 30:58]
  wire [31:0] inst_packet_6_inst_addr = {inst_packet_0_inst_addr_hi_hi,3'h6,2'h0}; // @[Cat.scala 30:58]
  wire [31:0] inst_packet_7_inst_addr = {inst_packet_0_inst_addr_hi_hi,3'h7,2'h0}; // @[Cat.scala 30:58]
  wire  _GEN_0 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_0 & tail[0] ? io_bpu_inst_packet_i_bits_predict_mask_0 :
    fetch_buffer_0_predict_taken; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25 FetchBuffer.scala 50:25]
  wire [3:0] _GEN_4 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_0 & tail[0] ? io_bpu_inst_packet_i_bits_gh_backup :
    fetch_buffer_0_gh_backup; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25 FetchBuffer.scala 50:25]
  wire [31:0] _GEN_5 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_0 & tail[0] ? inst_packet_0_inst_addr :
    fetch_buffer_0_inst_addr; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25 FetchBuffer.scala 50:25]
  wire [31:0] _GEN_6 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_0 & tail[0] ? io_bpu_inst_packet_i_bits_data_0 :
    fetch_buffer_0_inst; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25 FetchBuffer.scala 50:25]
  wire  _GEN_7 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_0 & tail[1] ? io_bpu_inst_packet_i_bits_predict_mask_0 :
    fetch_buffer_1_predict_taken; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25 FetchBuffer.scala 50:25]
  wire [3:0] _GEN_11 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_0 & tail[1] ? io_bpu_inst_packet_i_bits_gh_backup
     : fetch_buffer_1_gh_backup; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25 FetchBuffer.scala 50:25]
  wire [31:0] _GEN_12 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_0 & tail[1] ? inst_packet_0_inst_addr :
    fetch_buffer_1_inst_addr; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25 FetchBuffer.scala 50:25]
  wire [31:0] _GEN_13 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_0 & tail[1] ? io_bpu_inst_packet_i_bits_data_0 :
    fetch_buffer_1_inst; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25 FetchBuffer.scala 50:25]
  wire  _GEN_14 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_0 & tail[2] ? io_bpu_inst_packet_i_bits_predict_mask_0
     : fetch_buffer_2_predict_taken; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25 FetchBuffer.scala 50:25]
  wire [3:0] _GEN_18 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_0 & tail[2] ? io_bpu_inst_packet_i_bits_gh_backup
     : fetch_buffer_2_gh_backup; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25 FetchBuffer.scala 50:25]
  wire [31:0] _GEN_19 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_0 & tail[2] ? inst_packet_0_inst_addr :
    fetch_buffer_2_inst_addr; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25 FetchBuffer.scala 50:25]
  wire [31:0] _GEN_20 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_0 & tail[2] ? io_bpu_inst_packet_i_bits_data_0 :
    fetch_buffer_2_inst; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25 FetchBuffer.scala 50:25]
  wire  _GEN_21 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_0 & tail[3] ? io_bpu_inst_packet_i_bits_predict_mask_0
     : fetch_buffer_3_predict_taken; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25 FetchBuffer.scala 50:25]
  wire [3:0] _GEN_25 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_0 & tail[3] ? io_bpu_inst_packet_i_bits_gh_backup
     : fetch_buffer_3_gh_backup; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25 FetchBuffer.scala 50:25]
  wire [31:0] _GEN_26 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_0 & tail[3] ? inst_packet_0_inst_addr :
    fetch_buffer_3_inst_addr; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25 FetchBuffer.scala 50:25]
  wire [31:0] _GEN_27 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_0 & tail[3] ? io_bpu_inst_packet_i_bits_data_0 :
    fetch_buffer_3_inst; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25 FetchBuffer.scala 50:25]
  wire  _GEN_28 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_0 & tail[4] ? io_bpu_inst_packet_i_bits_predict_mask_0
     : fetch_buffer_4_predict_taken; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25 FetchBuffer.scala 50:25]
  wire [3:0] _GEN_32 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_0 & tail[4] ? io_bpu_inst_packet_i_bits_gh_backup
     : fetch_buffer_4_gh_backup; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25 FetchBuffer.scala 50:25]
  wire [31:0] _GEN_33 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_0 & tail[4] ? inst_packet_0_inst_addr :
    fetch_buffer_4_inst_addr; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25 FetchBuffer.scala 50:25]
  wire [31:0] _GEN_34 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_0 & tail[4] ? io_bpu_inst_packet_i_bits_data_0 :
    fetch_buffer_4_inst; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25 FetchBuffer.scala 50:25]
  wire  _GEN_35 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_0 & tail[5] ? io_bpu_inst_packet_i_bits_predict_mask_0
     : fetch_buffer_5_predict_taken; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25 FetchBuffer.scala 50:25]
  wire [3:0] _GEN_39 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_0 & tail[5] ? io_bpu_inst_packet_i_bits_gh_backup
     : fetch_buffer_5_gh_backup; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25 FetchBuffer.scala 50:25]
  wire [31:0] _GEN_40 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_0 & tail[5] ? inst_packet_0_inst_addr :
    fetch_buffer_5_inst_addr; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25 FetchBuffer.scala 50:25]
  wire [31:0] _GEN_41 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_0 & tail[5] ? io_bpu_inst_packet_i_bits_data_0 :
    fetch_buffer_5_inst; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25 FetchBuffer.scala 50:25]
  wire  _GEN_42 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_0 & tail[6] ? io_bpu_inst_packet_i_bits_predict_mask_0
     : fetch_buffer_6_predict_taken; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25 FetchBuffer.scala 50:25]
  wire [3:0] _GEN_46 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_0 & tail[6] ? io_bpu_inst_packet_i_bits_gh_backup
     : fetch_buffer_6_gh_backup; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25 FetchBuffer.scala 50:25]
  wire [31:0] _GEN_47 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_0 & tail[6] ? inst_packet_0_inst_addr :
    fetch_buffer_6_inst_addr; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25 FetchBuffer.scala 50:25]
  wire [31:0] _GEN_48 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_0 & tail[6] ? io_bpu_inst_packet_i_bits_data_0 :
    fetch_buffer_6_inst; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25 FetchBuffer.scala 50:25]
  wire  _GEN_49 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_0 & tail[7] ? io_bpu_inst_packet_i_bits_predict_mask_0
     : fetch_buffer_7_predict_taken; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25 FetchBuffer.scala 50:25]
  wire [3:0] _GEN_53 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_0 & tail[7] ? io_bpu_inst_packet_i_bits_gh_backup
     : fetch_buffer_7_gh_backup; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25 FetchBuffer.scala 50:25]
  wire [31:0] _GEN_54 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_0 & tail[7] ? inst_packet_0_inst_addr :
    fetch_buffer_7_inst_addr; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25 FetchBuffer.scala 50:25]
  wire [31:0] _GEN_55 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_0 & tail[7] ? io_bpu_inst_packet_i_bits_data_0 :
    fetch_buffer_7_inst; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25 FetchBuffer.scala 50:25]
  wire  _GEN_56 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_0 & tail[8] ? io_bpu_inst_packet_i_bits_predict_mask_0
     : fetch_buffer_8_predict_taken; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25 FetchBuffer.scala 50:25]
  wire [3:0] _GEN_60 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_0 & tail[8] ? io_bpu_inst_packet_i_bits_gh_backup
     : fetch_buffer_8_gh_backup; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25 FetchBuffer.scala 50:25]
  wire [31:0] _GEN_61 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_0 & tail[8] ? inst_packet_0_inst_addr :
    fetch_buffer_8_inst_addr; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25 FetchBuffer.scala 50:25]
  wire [31:0] _GEN_62 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_0 & tail[8] ? io_bpu_inst_packet_i_bits_data_0 :
    fetch_buffer_8_inst; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25 FetchBuffer.scala 50:25]
  wire  _GEN_63 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_0 & tail[9] ? io_bpu_inst_packet_i_bits_predict_mask_0
     : fetch_buffer_9_predict_taken; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25 FetchBuffer.scala 50:25]
  wire [3:0] _GEN_67 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_0 & tail[9] ? io_bpu_inst_packet_i_bits_gh_backup
     : fetch_buffer_9_gh_backup; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25 FetchBuffer.scala 50:25]
  wire [31:0] _GEN_68 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_0 & tail[9] ? inst_packet_0_inst_addr :
    fetch_buffer_9_inst_addr; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25 FetchBuffer.scala 50:25]
  wire [31:0] _GEN_69 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_0 & tail[9] ? io_bpu_inst_packet_i_bits_data_0 :
    fetch_buffer_9_inst; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25 FetchBuffer.scala 50:25]
  wire  _GEN_70 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_0 & tail[10] ? io_bpu_inst_packet_i_bits_predict_mask_0
     : fetch_buffer_10_predict_taken; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25 FetchBuffer.scala 50:25]
  wire [3:0] _GEN_74 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_0 & tail[10] ? io_bpu_inst_packet_i_bits_gh_backup
     : fetch_buffer_10_gh_backup; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25 FetchBuffer.scala 50:25]
  wire [31:0] _GEN_75 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_0 & tail[10] ? inst_packet_0_inst_addr :
    fetch_buffer_10_inst_addr; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25 FetchBuffer.scala 50:25]
  wire [31:0] _GEN_76 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_0 & tail[10] ? io_bpu_inst_packet_i_bits_data_0 :
    fetch_buffer_10_inst; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25 FetchBuffer.scala 50:25]
  wire  _GEN_77 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_0 & tail[11] ? io_bpu_inst_packet_i_bits_predict_mask_0
     : fetch_buffer_11_predict_taken; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25 FetchBuffer.scala 50:25]
  wire [3:0] _GEN_81 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_0 & tail[11] ? io_bpu_inst_packet_i_bits_gh_backup
     : fetch_buffer_11_gh_backup; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25 FetchBuffer.scala 50:25]
  wire [31:0] _GEN_82 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_0 & tail[11] ? inst_packet_0_inst_addr :
    fetch_buffer_11_inst_addr; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25 FetchBuffer.scala 50:25]
  wire [31:0] _GEN_83 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_0 & tail[11] ? io_bpu_inst_packet_i_bits_data_0 :
    fetch_buffer_11_inst; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25 FetchBuffer.scala 50:25]
  wire  _GEN_84 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_0 & tail[12] ? io_bpu_inst_packet_i_bits_predict_mask_0
     : fetch_buffer_12_predict_taken; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25 FetchBuffer.scala 50:25]
  wire [3:0] _GEN_88 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_0 & tail[12] ? io_bpu_inst_packet_i_bits_gh_backup
     : fetch_buffer_12_gh_backup; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25 FetchBuffer.scala 50:25]
  wire [31:0] _GEN_89 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_0 & tail[12] ? inst_packet_0_inst_addr :
    fetch_buffer_12_inst_addr; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25 FetchBuffer.scala 50:25]
  wire [31:0] _GEN_90 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_0 & tail[12] ? io_bpu_inst_packet_i_bits_data_0 :
    fetch_buffer_12_inst; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25 FetchBuffer.scala 50:25]
  wire  _GEN_91 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_0 & tail[13] ? io_bpu_inst_packet_i_bits_predict_mask_0
     : fetch_buffer_13_predict_taken; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25 FetchBuffer.scala 50:25]
  wire [3:0] _GEN_95 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_0 & tail[13] ? io_bpu_inst_packet_i_bits_gh_backup
     : fetch_buffer_13_gh_backup; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25 FetchBuffer.scala 50:25]
  wire [31:0] _GEN_96 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_0 & tail[13] ? inst_packet_0_inst_addr :
    fetch_buffer_13_inst_addr; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25 FetchBuffer.scala 50:25]
  wire [31:0] _GEN_97 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_0 & tail[13] ? io_bpu_inst_packet_i_bits_data_0 :
    fetch_buffer_13_inst; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25 FetchBuffer.scala 50:25]
  wire  _GEN_98 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_0 & tail[14] ? io_bpu_inst_packet_i_bits_predict_mask_0
     : fetch_buffer_14_predict_taken; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25 FetchBuffer.scala 50:25]
  wire [3:0] _GEN_102 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_0 & tail[14] ? io_bpu_inst_packet_i_bits_gh_backup
     : fetch_buffer_14_gh_backup; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25 FetchBuffer.scala 50:25]
  wire [31:0] _GEN_103 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_0 & tail[14] ? inst_packet_0_inst_addr :
    fetch_buffer_14_inst_addr; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25 FetchBuffer.scala 50:25]
  wire [31:0] _GEN_104 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_0 & tail[14] ? io_bpu_inst_packet_i_bits_data_0
     : fetch_buffer_14_inst; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25 FetchBuffer.scala 50:25]
  wire  _GEN_105 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_0 & tail[15] ? io_bpu_inst_packet_i_bits_predict_mask_0
     : fetch_buffer_15_predict_taken; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25 FetchBuffer.scala 50:25]
  wire [3:0] _GEN_109 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_0 & tail[15] ? io_bpu_inst_packet_i_bits_gh_backup
     : fetch_buffer_15_gh_backup; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25 FetchBuffer.scala 50:25]
  wire [31:0] _GEN_110 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_0 & tail[15] ? inst_packet_0_inst_addr :
    fetch_buffer_15_inst_addr; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25 FetchBuffer.scala 50:25]
  wire [31:0] _GEN_111 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_0 & tail[15] ? io_bpu_inst_packet_i_bits_data_0
     : fetch_buffer_15_inst; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25 FetchBuffer.scala 50:25]
  wire  _GEN_112 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_0 & lo ? io_bpu_inst_packet_i_bits_predict_mask_0 :
    fetch_buffer_16_predict_taken; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25 FetchBuffer.scala 50:25]
  wire [3:0] _GEN_116 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_0 & lo ? io_bpu_inst_packet_i_bits_gh_backup :
    fetch_buffer_16_gh_backup; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25 FetchBuffer.scala 50:25]
  wire [31:0] _GEN_117 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_0 & lo ? inst_packet_0_inst_addr :
    fetch_buffer_16_inst_addr; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25 FetchBuffer.scala 50:25]
  wire [31:0] _GEN_118 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_0 & lo ? io_bpu_inst_packet_i_bits_data_0 :
    fetch_buffer_16_inst; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25 FetchBuffer.scala 50:25]
  wire  _GEN_119 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_1 & enq_idxs_1[0] ?
    io_bpu_inst_packet_i_bits_predict_mask_1 : _GEN_0; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [3:0] _GEN_123 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_1 & enq_idxs_1[0] ?
    io_bpu_inst_packet_i_bits_gh_backup : _GEN_4; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_124 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_1 & enq_idxs_1[0] ? inst_packet_1_inst_addr :
    _GEN_5; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_125 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_1 & enq_idxs_1[0] ?
    io_bpu_inst_packet_i_bits_data_1 : _GEN_6; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire  _GEN_126 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_1 & enq_idxs_1[1] ?
    io_bpu_inst_packet_i_bits_predict_mask_1 : _GEN_7; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [3:0] _GEN_130 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_1 & enq_idxs_1[1] ?
    io_bpu_inst_packet_i_bits_gh_backup : _GEN_11; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_131 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_1 & enq_idxs_1[1] ? inst_packet_1_inst_addr :
    _GEN_12; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_132 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_1 & enq_idxs_1[1] ?
    io_bpu_inst_packet_i_bits_data_1 : _GEN_13; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire  _GEN_133 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_1 & enq_idxs_1[2] ?
    io_bpu_inst_packet_i_bits_predict_mask_1 : _GEN_14; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [3:0] _GEN_137 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_1 & enq_idxs_1[2] ?
    io_bpu_inst_packet_i_bits_gh_backup : _GEN_18; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_138 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_1 & enq_idxs_1[2] ? inst_packet_1_inst_addr :
    _GEN_19; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_139 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_1 & enq_idxs_1[2] ?
    io_bpu_inst_packet_i_bits_data_1 : _GEN_20; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire  _GEN_140 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_1 & enq_idxs_1[3] ?
    io_bpu_inst_packet_i_bits_predict_mask_1 : _GEN_21; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [3:0] _GEN_144 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_1 & enq_idxs_1[3] ?
    io_bpu_inst_packet_i_bits_gh_backup : _GEN_25; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_145 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_1 & enq_idxs_1[3] ? inst_packet_1_inst_addr :
    _GEN_26; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_146 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_1 & enq_idxs_1[3] ?
    io_bpu_inst_packet_i_bits_data_1 : _GEN_27; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire  _GEN_147 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_1 & enq_idxs_1[4] ?
    io_bpu_inst_packet_i_bits_predict_mask_1 : _GEN_28; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [3:0] _GEN_151 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_1 & enq_idxs_1[4] ?
    io_bpu_inst_packet_i_bits_gh_backup : _GEN_32; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_152 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_1 & enq_idxs_1[4] ? inst_packet_1_inst_addr :
    _GEN_33; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_153 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_1 & enq_idxs_1[4] ?
    io_bpu_inst_packet_i_bits_data_1 : _GEN_34; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire  _GEN_154 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_1 & enq_idxs_1[5] ?
    io_bpu_inst_packet_i_bits_predict_mask_1 : _GEN_35; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [3:0] _GEN_158 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_1 & enq_idxs_1[5] ?
    io_bpu_inst_packet_i_bits_gh_backup : _GEN_39; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_159 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_1 & enq_idxs_1[5] ? inst_packet_1_inst_addr :
    _GEN_40; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_160 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_1 & enq_idxs_1[5] ?
    io_bpu_inst_packet_i_bits_data_1 : _GEN_41; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire  _GEN_161 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_1 & enq_idxs_1[6] ?
    io_bpu_inst_packet_i_bits_predict_mask_1 : _GEN_42; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [3:0] _GEN_165 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_1 & enq_idxs_1[6] ?
    io_bpu_inst_packet_i_bits_gh_backup : _GEN_46; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_166 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_1 & enq_idxs_1[6] ? inst_packet_1_inst_addr :
    _GEN_47; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_167 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_1 & enq_idxs_1[6] ?
    io_bpu_inst_packet_i_bits_data_1 : _GEN_48; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire  _GEN_168 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_1 & enq_idxs_1[7] ?
    io_bpu_inst_packet_i_bits_predict_mask_1 : _GEN_49; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [3:0] _GEN_172 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_1 & enq_idxs_1[7] ?
    io_bpu_inst_packet_i_bits_gh_backup : _GEN_53; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_173 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_1 & enq_idxs_1[7] ? inst_packet_1_inst_addr :
    _GEN_54; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_174 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_1 & enq_idxs_1[7] ?
    io_bpu_inst_packet_i_bits_data_1 : _GEN_55; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire  _GEN_175 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_1 & enq_idxs_1[8] ?
    io_bpu_inst_packet_i_bits_predict_mask_1 : _GEN_56; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [3:0] _GEN_179 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_1 & enq_idxs_1[8] ?
    io_bpu_inst_packet_i_bits_gh_backup : _GEN_60; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_180 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_1 & enq_idxs_1[8] ? inst_packet_1_inst_addr :
    _GEN_61; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_181 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_1 & enq_idxs_1[8] ?
    io_bpu_inst_packet_i_bits_data_1 : _GEN_62; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire  _GEN_182 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_1 & enq_idxs_1[9] ?
    io_bpu_inst_packet_i_bits_predict_mask_1 : _GEN_63; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [3:0] _GEN_186 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_1 & enq_idxs_1[9] ?
    io_bpu_inst_packet_i_bits_gh_backup : _GEN_67; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_187 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_1 & enq_idxs_1[9] ? inst_packet_1_inst_addr :
    _GEN_68; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_188 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_1 & enq_idxs_1[9] ?
    io_bpu_inst_packet_i_bits_data_1 : _GEN_69; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire  _GEN_189 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_1 & enq_idxs_1[10] ?
    io_bpu_inst_packet_i_bits_predict_mask_1 : _GEN_70; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [3:0] _GEN_193 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_1 & enq_idxs_1[10] ?
    io_bpu_inst_packet_i_bits_gh_backup : _GEN_74; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_194 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_1 & enq_idxs_1[10] ? inst_packet_1_inst_addr :
    _GEN_75; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_195 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_1 & enq_idxs_1[10] ?
    io_bpu_inst_packet_i_bits_data_1 : _GEN_76; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire  _GEN_196 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_1 & enq_idxs_1[11] ?
    io_bpu_inst_packet_i_bits_predict_mask_1 : _GEN_77; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [3:0] _GEN_200 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_1 & enq_idxs_1[11] ?
    io_bpu_inst_packet_i_bits_gh_backup : _GEN_81; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_201 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_1 & enq_idxs_1[11] ? inst_packet_1_inst_addr :
    _GEN_82; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_202 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_1 & enq_idxs_1[11] ?
    io_bpu_inst_packet_i_bits_data_1 : _GEN_83; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire  _GEN_203 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_1 & enq_idxs_1[12] ?
    io_bpu_inst_packet_i_bits_predict_mask_1 : _GEN_84; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [3:0] _GEN_207 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_1 & enq_idxs_1[12] ?
    io_bpu_inst_packet_i_bits_gh_backup : _GEN_88; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_208 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_1 & enq_idxs_1[12] ? inst_packet_1_inst_addr :
    _GEN_89; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_209 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_1 & enq_idxs_1[12] ?
    io_bpu_inst_packet_i_bits_data_1 : _GEN_90; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire  _GEN_210 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_1 & enq_idxs_1[13] ?
    io_bpu_inst_packet_i_bits_predict_mask_1 : _GEN_91; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [3:0] _GEN_214 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_1 & enq_idxs_1[13] ?
    io_bpu_inst_packet_i_bits_gh_backup : _GEN_95; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_215 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_1 & enq_idxs_1[13] ? inst_packet_1_inst_addr :
    _GEN_96; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_216 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_1 & enq_idxs_1[13] ?
    io_bpu_inst_packet_i_bits_data_1 : _GEN_97; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire  _GEN_217 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_1 & enq_idxs_1[14] ?
    io_bpu_inst_packet_i_bits_predict_mask_1 : _GEN_98; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [3:0] _GEN_221 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_1 & enq_idxs_1[14] ?
    io_bpu_inst_packet_i_bits_gh_backup : _GEN_102; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_222 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_1 & enq_idxs_1[14] ? inst_packet_1_inst_addr :
    _GEN_103; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_223 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_1 & enq_idxs_1[14] ?
    io_bpu_inst_packet_i_bits_data_1 : _GEN_104; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire  _GEN_224 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_1 & enq_idxs_1[15] ?
    io_bpu_inst_packet_i_bits_predict_mask_1 : _GEN_105; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [3:0] _GEN_228 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_1 & enq_idxs_1[15] ?
    io_bpu_inst_packet_i_bits_gh_backup : _GEN_109; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_229 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_1 & enq_idxs_1[15] ? inst_packet_1_inst_addr :
    _GEN_110; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_230 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_1 & enq_idxs_1[15] ?
    io_bpu_inst_packet_i_bits_data_1 : _GEN_111; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire  _GEN_231 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_1 & lo_1 ? io_bpu_inst_packet_i_bits_predict_mask_1 :
    _GEN_112; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [3:0] _GEN_235 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_1 & lo_1 ? io_bpu_inst_packet_i_bits_gh_backup :
    _GEN_116; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_236 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_1 & lo_1 ? inst_packet_1_inst_addr : _GEN_117; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_237 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_1 & lo_1 ? io_bpu_inst_packet_i_bits_data_1 :
    _GEN_118; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire  _GEN_238 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_2 & enq_idxs_2[0] ?
    io_bpu_inst_packet_i_bits_predict_mask_2 : _GEN_119; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [3:0] _GEN_242 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_2 & enq_idxs_2[0] ?
    io_bpu_inst_packet_i_bits_gh_backup : _GEN_123; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_243 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_2 & enq_idxs_2[0] ? inst_packet_2_inst_addr :
    _GEN_124; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_244 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_2 & enq_idxs_2[0] ?
    io_bpu_inst_packet_i_bits_data_2 : _GEN_125; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire  _GEN_245 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_2 & enq_idxs_2[1] ?
    io_bpu_inst_packet_i_bits_predict_mask_2 : _GEN_126; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [3:0] _GEN_249 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_2 & enq_idxs_2[1] ?
    io_bpu_inst_packet_i_bits_gh_backup : _GEN_130; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_250 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_2 & enq_idxs_2[1] ? inst_packet_2_inst_addr :
    _GEN_131; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_251 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_2 & enq_idxs_2[1] ?
    io_bpu_inst_packet_i_bits_data_2 : _GEN_132; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire  _GEN_252 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_2 & enq_idxs_2[2] ?
    io_bpu_inst_packet_i_bits_predict_mask_2 : _GEN_133; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [3:0] _GEN_256 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_2 & enq_idxs_2[2] ?
    io_bpu_inst_packet_i_bits_gh_backup : _GEN_137; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_257 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_2 & enq_idxs_2[2] ? inst_packet_2_inst_addr :
    _GEN_138; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_258 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_2 & enq_idxs_2[2] ?
    io_bpu_inst_packet_i_bits_data_2 : _GEN_139; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire  _GEN_259 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_2 & enq_idxs_2[3] ?
    io_bpu_inst_packet_i_bits_predict_mask_2 : _GEN_140; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [3:0] _GEN_263 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_2 & enq_idxs_2[3] ?
    io_bpu_inst_packet_i_bits_gh_backup : _GEN_144; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_264 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_2 & enq_idxs_2[3] ? inst_packet_2_inst_addr :
    _GEN_145; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_265 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_2 & enq_idxs_2[3] ?
    io_bpu_inst_packet_i_bits_data_2 : _GEN_146; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire  _GEN_266 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_2 & enq_idxs_2[4] ?
    io_bpu_inst_packet_i_bits_predict_mask_2 : _GEN_147; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [3:0] _GEN_270 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_2 & enq_idxs_2[4] ?
    io_bpu_inst_packet_i_bits_gh_backup : _GEN_151; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_271 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_2 & enq_idxs_2[4] ? inst_packet_2_inst_addr :
    _GEN_152; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_272 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_2 & enq_idxs_2[4] ?
    io_bpu_inst_packet_i_bits_data_2 : _GEN_153; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire  _GEN_273 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_2 & enq_idxs_2[5] ?
    io_bpu_inst_packet_i_bits_predict_mask_2 : _GEN_154; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [3:0] _GEN_277 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_2 & enq_idxs_2[5] ?
    io_bpu_inst_packet_i_bits_gh_backup : _GEN_158; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_278 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_2 & enq_idxs_2[5] ? inst_packet_2_inst_addr :
    _GEN_159; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_279 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_2 & enq_idxs_2[5] ?
    io_bpu_inst_packet_i_bits_data_2 : _GEN_160; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire  _GEN_280 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_2 & enq_idxs_2[6] ?
    io_bpu_inst_packet_i_bits_predict_mask_2 : _GEN_161; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [3:0] _GEN_284 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_2 & enq_idxs_2[6] ?
    io_bpu_inst_packet_i_bits_gh_backup : _GEN_165; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_285 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_2 & enq_idxs_2[6] ? inst_packet_2_inst_addr :
    _GEN_166; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_286 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_2 & enq_idxs_2[6] ?
    io_bpu_inst_packet_i_bits_data_2 : _GEN_167; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire  _GEN_287 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_2 & enq_idxs_2[7] ?
    io_bpu_inst_packet_i_bits_predict_mask_2 : _GEN_168; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [3:0] _GEN_291 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_2 & enq_idxs_2[7] ?
    io_bpu_inst_packet_i_bits_gh_backup : _GEN_172; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_292 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_2 & enq_idxs_2[7] ? inst_packet_2_inst_addr :
    _GEN_173; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_293 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_2 & enq_idxs_2[7] ?
    io_bpu_inst_packet_i_bits_data_2 : _GEN_174; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire  _GEN_294 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_2 & enq_idxs_2[8] ?
    io_bpu_inst_packet_i_bits_predict_mask_2 : _GEN_175; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [3:0] _GEN_298 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_2 & enq_idxs_2[8] ?
    io_bpu_inst_packet_i_bits_gh_backup : _GEN_179; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_299 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_2 & enq_idxs_2[8] ? inst_packet_2_inst_addr :
    _GEN_180; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_300 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_2 & enq_idxs_2[8] ?
    io_bpu_inst_packet_i_bits_data_2 : _GEN_181; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire  _GEN_301 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_2 & enq_idxs_2[9] ?
    io_bpu_inst_packet_i_bits_predict_mask_2 : _GEN_182; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [3:0] _GEN_305 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_2 & enq_idxs_2[9] ?
    io_bpu_inst_packet_i_bits_gh_backup : _GEN_186; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_306 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_2 & enq_idxs_2[9] ? inst_packet_2_inst_addr :
    _GEN_187; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_307 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_2 & enq_idxs_2[9] ?
    io_bpu_inst_packet_i_bits_data_2 : _GEN_188; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire  _GEN_308 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_2 & enq_idxs_2[10] ?
    io_bpu_inst_packet_i_bits_predict_mask_2 : _GEN_189; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [3:0] _GEN_312 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_2 & enq_idxs_2[10] ?
    io_bpu_inst_packet_i_bits_gh_backup : _GEN_193; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_313 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_2 & enq_idxs_2[10] ? inst_packet_2_inst_addr :
    _GEN_194; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_314 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_2 & enq_idxs_2[10] ?
    io_bpu_inst_packet_i_bits_data_2 : _GEN_195; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire  _GEN_315 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_2 & enq_idxs_2[11] ?
    io_bpu_inst_packet_i_bits_predict_mask_2 : _GEN_196; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [3:0] _GEN_319 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_2 & enq_idxs_2[11] ?
    io_bpu_inst_packet_i_bits_gh_backup : _GEN_200; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_320 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_2 & enq_idxs_2[11] ? inst_packet_2_inst_addr :
    _GEN_201; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_321 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_2 & enq_idxs_2[11] ?
    io_bpu_inst_packet_i_bits_data_2 : _GEN_202; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire  _GEN_322 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_2 & enq_idxs_2[12] ?
    io_bpu_inst_packet_i_bits_predict_mask_2 : _GEN_203; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [3:0] _GEN_326 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_2 & enq_idxs_2[12] ?
    io_bpu_inst_packet_i_bits_gh_backup : _GEN_207; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_327 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_2 & enq_idxs_2[12] ? inst_packet_2_inst_addr :
    _GEN_208; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_328 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_2 & enq_idxs_2[12] ?
    io_bpu_inst_packet_i_bits_data_2 : _GEN_209; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire  _GEN_329 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_2 & enq_idxs_2[13] ?
    io_bpu_inst_packet_i_bits_predict_mask_2 : _GEN_210; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [3:0] _GEN_333 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_2 & enq_idxs_2[13] ?
    io_bpu_inst_packet_i_bits_gh_backup : _GEN_214; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_334 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_2 & enq_idxs_2[13] ? inst_packet_2_inst_addr :
    _GEN_215; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_335 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_2 & enq_idxs_2[13] ?
    io_bpu_inst_packet_i_bits_data_2 : _GEN_216; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire  _GEN_336 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_2 & enq_idxs_2[14] ?
    io_bpu_inst_packet_i_bits_predict_mask_2 : _GEN_217; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [3:0] _GEN_340 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_2 & enq_idxs_2[14] ?
    io_bpu_inst_packet_i_bits_gh_backup : _GEN_221; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_341 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_2 & enq_idxs_2[14] ? inst_packet_2_inst_addr :
    _GEN_222; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_342 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_2 & enq_idxs_2[14] ?
    io_bpu_inst_packet_i_bits_data_2 : _GEN_223; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire  _GEN_343 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_2 & enq_idxs_2[15] ?
    io_bpu_inst_packet_i_bits_predict_mask_2 : _GEN_224; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [3:0] _GEN_347 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_2 & enq_idxs_2[15] ?
    io_bpu_inst_packet_i_bits_gh_backup : _GEN_228; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_348 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_2 & enq_idxs_2[15] ? inst_packet_2_inst_addr :
    _GEN_229; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_349 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_2 & enq_idxs_2[15] ?
    io_bpu_inst_packet_i_bits_data_2 : _GEN_230; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire  _GEN_350 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_2 & lo_2 ? io_bpu_inst_packet_i_bits_predict_mask_2 :
    _GEN_231; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [3:0] _GEN_354 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_2 & lo_2 ? io_bpu_inst_packet_i_bits_gh_backup :
    _GEN_235; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_355 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_2 & lo_2 ? inst_packet_2_inst_addr : _GEN_236; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_356 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_2 & lo_2 ? io_bpu_inst_packet_i_bits_data_2 :
    _GEN_237; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire  _GEN_357 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_3 & enq_idxs_3[0] ?
    io_bpu_inst_packet_i_bits_predict_mask_3 : _GEN_238; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [3:0] _GEN_361 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_3 & enq_idxs_3[0] ?
    io_bpu_inst_packet_i_bits_gh_backup : _GEN_242; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_362 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_3 & enq_idxs_3[0] ? inst_packet_3_inst_addr :
    _GEN_243; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_363 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_3 & enq_idxs_3[0] ?
    io_bpu_inst_packet_i_bits_data_3 : _GEN_244; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire  _GEN_364 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_3 & enq_idxs_3[1] ?
    io_bpu_inst_packet_i_bits_predict_mask_3 : _GEN_245; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [3:0] _GEN_368 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_3 & enq_idxs_3[1] ?
    io_bpu_inst_packet_i_bits_gh_backup : _GEN_249; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_369 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_3 & enq_idxs_3[1] ? inst_packet_3_inst_addr :
    _GEN_250; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_370 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_3 & enq_idxs_3[1] ?
    io_bpu_inst_packet_i_bits_data_3 : _GEN_251; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire  _GEN_371 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_3 & enq_idxs_3[2] ?
    io_bpu_inst_packet_i_bits_predict_mask_3 : _GEN_252; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [3:0] _GEN_375 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_3 & enq_idxs_3[2] ?
    io_bpu_inst_packet_i_bits_gh_backup : _GEN_256; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_376 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_3 & enq_idxs_3[2] ? inst_packet_3_inst_addr :
    _GEN_257; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_377 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_3 & enq_idxs_3[2] ?
    io_bpu_inst_packet_i_bits_data_3 : _GEN_258; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire  _GEN_378 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_3 & enq_idxs_3[3] ?
    io_bpu_inst_packet_i_bits_predict_mask_3 : _GEN_259; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [3:0] _GEN_382 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_3 & enq_idxs_3[3] ?
    io_bpu_inst_packet_i_bits_gh_backup : _GEN_263; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_383 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_3 & enq_idxs_3[3] ? inst_packet_3_inst_addr :
    _GEN_264; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_384 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_3 & enq_idxs_3[3] ?
    io_bpu_inst_packet_i_bits_data_3 : _GEN_265; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire  _GEN_385 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_3 & enq_idxs_3[4] ?
    io_bpu_inst_packet_i_bits_predict_mask_3 : _GEN_266; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [3:0] _GEN_389 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_3 & enq_idxs_3[4] ?
    io_bpu_inst_packet_i_bits_gh_backup : _GEN_270; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_390 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_3 & enq_idxs_3[4] ? inst_packet_3_inst_addr :
    _GEN_271; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_391 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_3 & enq_idxs_3[4] ?
    io_bpu_inst_packet_i_bits_data_3 : _GEN_272; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire  _GEN_392 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_3 & enq_idxs_3[5] ?
    io_bpu_inst_packet_i_bits_predict_mask_3 : _GEN_273; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [3:0] _GEN_396 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_3 & enq_idxs_3[5] ?
    io_bpu_inst_packet_i_bits_gh_backup : _GEN_277; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_397 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_3 & enq_idxs_3[5] ? inst_packet_3_inst_addr :
    _GEN_278; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_398 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_3 & enq_idxs_3[5] ?
    io_bpu_inst_packet_i_bits_data_3 : _GEN_279; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire  _GEN_399 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_3 & enq_idxs_3[6] ?
    io_bpu_inst_packet_i_bits_predict_mask_3 : _GEN_280; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [3:0] _GEN_403 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_3 & enq_idxs_3[6] ?
    io_bpu_inst_packet_i_bits_gh_backup : _GEN_284; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_404 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_3 & enq_idxs_3[6] ? inst_packet_3_inst_addr :
    _GEN_285; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_405 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_3 & enq_idxs_3[6] ?
    io_bpu_inst_packet_i_bits_data_3 : _GEN_286; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire  _GEN_406 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_3 & enq_idxs_3[7] ?
    io_bpu_inst_packet_i_bits_predict_mask_3 : _GEN_287; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [3:0] _GEN_410 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_3 & enq_idxs_3[7] ?
    io_bpu_inst_packet_i_bits_gh_backup : _GEN_291; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_411 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_3 & enq_idxs_3[7] ? inst_packet_3_inst_addr :
    _GEN_292; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_412 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_3 & enq_idxs_3[7] ?
    io_bpu_inst_packet_i_bits_data_3 : _GEN_293; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire  _GEN_413 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_3 & enq_idxs_3[8] ?
    io_bpu_inst_packet_i_bits_predict_mask_3 : _GEN_294; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [3:0] _GEN_417 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_3 & enq_idxs_3[8] ?
    io_bpu_inst_packet_i_bits_gh_backup : _GEN_298; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_418 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_3 & enq_idxs_3[8] ? inst_packet_3_inst_addr :
    _GEN_299; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_419 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_3 & enq_idxs_3[8] ?
    io_bpu_inst_packet_i_bits_data_3 : _GEN_300; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire  _GEN_420 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_3 & enq_idxs_3[9] ?
    io_bpu_inst_packet_i_bits_predict_mask_3 : _GEN_301; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [3:0] _GEN_424 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_3 & enq_idxs_3[9] ?
    io_bpu_inst_packet_i_bits_gh_backup : _GEN_305; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_425 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_3 & enq_idxs_3[9] ? inst_packet_3_inst_addr :
    _GEN_306; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_426 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_3 & enq_idxs_3[9] ?
    io_bpu_inst_packet_i_bits_data_3 : _GEN_307; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire  _GEN_427 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_3 & enq_idxs_3[10] ?
    io_bpu_inst_packet_i_bits_predict_mask_3 : _GEN_308; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [3:0] _GEN_431 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_3 & enq_idxs_3[10] ?
    io_bpu_inst_packet_i_bits_gh_backup : _GEN_312; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_432 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_3 & enq_idxs_3[10] ? inst_packet_3_inst_addr :
    _GEN_313; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_433 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_3 & enq_idxs_3[10] ?
    io_bpu_inst_packet_i_bits_data_3 : _GEN_314; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire  _GEN_434 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_3 & enq_idxs_3[11] ?
    io_bpu_inst_packet_i_bits_predict_mask_3 : _GEN_315; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [3:0] _GEN_438 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_3 & enq_idxs_3[11] ?
    io_bpu_inst_packet_i_bits_gh_backup : _GEN_319; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_439 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_3 & enq_idxs_3[11] ? inst_packet_3_inst_addr :
    _GEN_320; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_440 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_3 & enq_idxs_3[11] ?
    io_bpu_inst_packet_i_bits_data_3 : _GEN_321; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire  _GEN_441 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_3 & enq_idxs_3[12] ?
    io_bpu_inst_packet_i_bits_predict_mask_3 : _GEN_322; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [3:0] _GEN_445 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_3 & enq_idxs_3[12] ?
    io_bpu_inst_packet_i_bits_gh_backup : _GEN_326; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_446 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_3 & enq_idxs_3[12] ? inst_packet_3_inst_addr :
    _GEN_327; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_447 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_3 & enq_idxs_3[12] ?
    io_bpu_inst_packet_i_bits_data_3 : _GEN_328; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire  _GEN_448 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_3 & enq_idxs_3[13] ?
    io_bpu_inst_packet_i_bits_predict_mask_3 : _GEN_329; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [3:0] _GEN_452 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_3 & enq_idxs_3[13] ?
    io_bpu_inst_packet_i_bits_gh_backup : _GEN_333; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_453 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_3 & enq_idxs_3[13] ? inst_packet_3_inst_addr :
    _GEN_334; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_454 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_3 & enq_idxs_3[13] ?
    io_bpu_inst_packet_i_bits_data_3 : _GEN_335; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire  _GEN_455 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_3 & enq_idxs_3[14] ?
    io_bpu_inst_packet_i_bits_predict_mask_3 : _GEN_336; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [3:0] _GEN_459 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_3 & enq_idxs_3[14] ?
    io_bpu_inst_packet_i_bits_gh_backup : _GEN_340; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_460 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_3 & enq_idxs_3[14] ? inst_packet_3_inst_addr :
    _GEN_341; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_461 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_3 & enq_idxs_3[14] ?
    io_bpu_inst_packet_i_bits_data_3 : _GEN_342; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire  _GEN_462 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_3 & enq_idxs_3[15] ?
    io_bpu_inst_packet_i_bits_predict_mask_3 : _GEN_343; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [3:0] _GEN_466 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_3 & enq_idxs_3[15] ?
    io_bpu_inst_packet_i_bits_gh_backup : _GEN_347; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_467 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_3 & enq_idxs_3[15] ? inst_packet_3_inst_addr :
    _GEN_348; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_468 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_3 & enq_idxs_3[15] ?
    io_bpu_inst_packet_i_bits_data_3 : _GEN_349; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire  _GEN_469 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_3 & lo_3 ? io_bpu_inst_packet_i_bits_predict_mask_3 :
    _GEN_350; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [3:0] _GEN_473 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_3 & lo_3 ? io_bpu_inst_packet_i_bits_gh_backup :
    _GEN_354; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_474 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_3 & lo_3 ? inst_packet_3_inst_addr : _GEN_355; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_475 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_3 & lo_3 ? io_bpu_inst_packet_i_bits_data_3 :
    _GEN_356; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [3:0] _GEN_480 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_4 & enq_idxs_4[0] ?
    io_bpu_inst_packet_i_bits_gh_backup : _GEN_361; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_481 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_4 & enq_idxs_4[0] ? inst_packet_4_inst_addr :
    _GEN_362; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_482 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_4 & enq_idxs_4[0] ?
    io_bpu_inst_packet_i_bits_data_4 : _GEN_363; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [3:0] _GEN_487 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_4 & enq_idxs_4[1] ?
    io_bpu_inst_packet_i_bits_gh_backup : _GEN_368; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_488 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_4 & enq_idxs_4[1] ? inst_packet_4_inst_addr :
    _GEN_369; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_489 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_4 & enq_idxs_4[1] ?
    io_bpu_inst_packet_i_bits_data_4 : _GEN_370; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [3:0] _GEN_494 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_4 & enq_idxs_4[2] ?
    io_bpu_inst_packet_i_bits_gh_backup : _GEN_375; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_495 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_4 & enq_idxs_4[2] ? inst_packet_4_inst_addr :
    _GEN_376; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_496 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_4 & enq_idxs_4[2] ?
    io_bpu_inst_packet_i_bits_data_4 : _GEN_377; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [3:0] _GEN_501 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_4 & enq_idxs_4[3] ?
    io_bpu_inst_packet_i_bits_gh_backup : _GEN_382; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_502 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_4 & enq_idxs_4[3] ? inst_packet_4_inst_addr :
    _GEN_383; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_503 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_4 & enq_idxs_4[3] ?
    io_bpu_inst_packet_i_bits_data_4 : _GEN_384; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [3:0] _GEN_508 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_4 & enq_idxs_4[4] ?
    io_bpu_inst_packet_i_bits_gh_backup : _GEN_389; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_509 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_4 & enq_idxs_4[4] ? inst_packet_4_inst_addr :
    _GEN_390; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_510 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_4 & enq_idxs_4[4] ?
    io_bpu_inst_packet_i_bits_data_4 : _GEN_391; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [3:0] _GEN_515 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_4 & enq_idxs_4[5] ?
    io_bpu_inst_packet_i_bits_gh_backup : _GEN_396; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_516 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_4 & enq_idxs_4[5] ? inst_packet_4_inst_addr :
    _GEN_397; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_517 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_4 & enq_idxs_4[5] ?
    io_bpu_inst_packet_i_bits_data_4 : _GEN_398; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [3:0] _GEN_522 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_4 & enq_idxs_4[6] ?
    io_bpu_inst_packet_i_bits_gh_backup : _GEN_403; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_523 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_4 & enq_idxs_4[6] ? inst_packet_4_inst_addr :
    _GEN_404; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_524 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_4 & enq_idxs_4[6] ?
    io_bpu_inst_packet_i_bits_data_4 : _GEN_405; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [3:0] _GEN_529 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_4 & enq_idxs_4[7] ?
    io_bpu_inst_packet_i_bits_gh_backup : _GEN_410; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_530 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_4 & enq_idxs_4[7] ? inst_packet_4_inst_addr :
    _GEN_411; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_531 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_4 & enq_idxs_4[7] ?
    io_bpu_inst_packet_i_bits_data_4 : _GEN_412; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [3:0] _GEN_536 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_4 & enq_idxs_4[8] ?
    io_bpu_inst_packet_i_bits_gh_backup : _GEN_417; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_537 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_4 & enq_idxs_4[8] ? inst_packet_4_inst_addr :
    _GEN_418; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_538 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_4 & enq_idxs_4[8] ?
    io_bpu_inst_packet_i_bits_data_4 : _GEN_419; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [3:0] _GEN_543 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_4 & enq_idxs_4[9] ?
    io_bpu_inst_packet_i_bits_gh_backup : _GEN_424; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_544 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_4 & enq_idxs_4[9] ? inst_packet_4_inst_addr :
    _GEN_425; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_545 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_4 & enq_idxs_4[9] ?
    io_bpu_inst_packet_i_bits_data_4 : _GEN_426; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [3:0] _GEN_550 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_4 & enq_idxs_4[10] ?
    io_bpu_inst_packet_i_bits_gh_backup : _GEN_431; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_551 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_4 & enq_idxs_4[10] ? inst_packet_4_inst_addr :
    _GEN_432; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_552 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_4 & enq_idxs_4[10] ?
    io_bpu_inst_packet_i_bits_data_4 : _GEN_433; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [3:0] _GEN_557 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_4 & enq_idxs_4[11] ?
    io_bpu_inst_packet_i_bits_gh_backup : _GEN_438; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_558 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_4 & enq_idxs_4[11] ? inst_packet_4_inst_addr :
    _GEN_439; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_559 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_4 & enq_idxs_4[11] ?
    io_bpu_inst_packet_i_bits_data_4 : _GEN_440; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [3:0] _GEN_564 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_4 & enq_idxs_4[12] ?
    io_bpu_inst_packet_i_bits_gh_backup : _GEN_445; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_565 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_4 & enq_idxs_4[12] ? inst_packet_4_inst_addr :
    _GEN_446; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_566 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_4 & enq_idxs_4[12] ?
    io_bpu_inst_packet_i_bits_data_4 : _GEN_447; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [3:0] _GEN_571 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_4 & enq_idxs_4[13] ?
    io_bpu_inst_packet_i_bits_gh_backup : _GEN_452; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_572 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_4 & enq_idxs_4[13] ? inst_packet_4_inst_addr :
    _GEN_453; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_573 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_4 & enq_idxs_4[13] ?
    io_bpu_inst_packet_i_bits_data_4 : _GEN_454; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [3:0] _GEN_578 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_4 & enq_idxs_4[14] ?
    io_bpu_inst_packet_i_bits_gh_backup : _GEN_459; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_579 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_4 & enq_idxs_4[14] ? inst_packet_4_inst_addr :
    _GEN_460; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_580 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_4 & enq_idxs_4[14] ?
    io_bpu_inst_packet_i_bits_data_4 : _GEN_461; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [3:0] _GEN_585 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_4 & enq_idxs_4[15] ?
    io_bpu_inst_packet_i_bits_gh_backup : _GEN_466; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_586 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_4 & enq_idxs_4[15] ? inst_packet_4_inst_addr :
    _GEN_467; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_587 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_4 & enq_idxs_4[15] ?
    io_bpu_inst_packet_i_bits_data_4 : _GEN_468; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [3:0] _GEN_592 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_4 & lo_4 ? io_bpu_inst_packet_i_bits_gh_backup :
    _GEN_473; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_593 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_4 & lo_4 ? inst_packet_4_inst_addr : _GEN_474; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [31:0] _GEN_594 = do_enq & io_bpu_inst_packet_i_bits_valid_mask_4 & lo_4 ? io_bpu_inst_packet_i_bits_data_4 :
    _GEN_475; // @[FetchBuffer.scala 84:65 FetchBuffer.scala 85:25]
  wire [15:0] deq_idxs_hi = deq_idxs_0[15:0]; // @[FetchBuffer.scala 42:12]
  wire  deq_idxs_lo = deq_idxs_0[16]; // @[FetchBuffer.scala 42:29]
  wire [16:0] deq_idxs_1 = {deq_idxs_hi,deq_idxs_lo}; // @[Cat.scala 30:58]
  wire  hit_tail_mask_0 = hit_head & ~is_full; // @[FetchBuffer.scala 97:47]
  wire  hit_tail_mask_1 = deq_idxs_1 == tail & ~is_full; // @[FetchBuffer.scala 97:47]
  wire  deq_invalid_1 = hit_tail_mask_0 | hit_tail_mask_1; // @[FetchBuffer.scala 98:57]
  wire  do_deq = io_fb_resp_deq_valid_0 | io_fb_resp_deq_valid_1; // @[FetchBuffer.scala 100:52]
  wire  _GEN_960 = deq_idxs_0[1] ? fetch_buffer_1_predict_taken : fetch_buffer_0_predict_taken; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire  _GEN_963 = deq_idxs_0[1] ? ~hit_tail_mask_0 : ~hit_tail_mask_0; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 105:44]
  wire [3:0] _GEN_964 = deq_idxs_0[1] ? fetch_buffer_1_gh_backup : fetch_buffer_0_gh_backup; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire [31:0] _GEN_965 = deq_idxs_0[1] ? fetch_buffer_1_inst_addr : fetch_buffer_0_inst_addr; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire [31:0] _GEN_966 = deq_idxs_0[1] ? fetch_buffer_1_inst : fetch_buffer_0_inst; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire  _GEN_967 = deq_idxs_0[2] ? fetch_buffer_2_predict_taken : _GEN_960; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire  _GEN_970 = deq_idxs_0[2] ? ~hit_tail_mask_0 : _GEN_963; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 105:44]
  wire [3:0] _GEN_971 = deq_idxs_0[2] ? fetch_buffer_2_gh_backup : _GEN_964; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire [31:0] _GEN_972 = deq_idxs_0[2] ? fetch_buffer_2_inst_addr : _GEN_965; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire [31:0] _GEN_973 = deq_idxs_0[2] ? fetch_buffer_2_inst : _GEN_966; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire  _GEN_974 = deq_idxs_0[3] ? fetch_buffer_3_predict_taken : _GEN_967; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire  _GEN_977 = deq_idxs_0[3] ? ~hit_tail_mask_0 : _GEN_970; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 105:44]
  wire [3:0] _GEN_978 = deq_idxs_0[3] ? fetch_buffer_3_gh_backup : _GEN_971; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire [31:0] _GEN_979 = deq_idxs_0[3] ? fetch_buffer_3_inst_addr : _GEN_972; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire [31:0] _GEN_980 = deq_idxs_0[3] ? fetch_buffer_3_inst : _GEN_973; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire  _GEN_981 = deq_idxs_0[4] ? fetch_buffer_4_predict_taken : _GEN_974; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire  _GEN_984 = deq_idxs_0[4] ? ~hit_tail_mask_0 : _GEN_977; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 105:44]
  wire [3:0] _GEN_985 = deq_idxs_0[4] ? fetch_buffer_4_gh_backup : _GEN_978; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire [31:0] _GEN_986 = deq_idxs_0[4] ? fetch_buffer_4_inst_addr : _GEN_979; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire [31:0] _GEN_987 = deq_idxs_0[4] ? fetch_buffer_4_inst : _GEN_980; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire  _GEN_988 = deq_idxs_0[5] ? fetch_buffer_5_predict_taken : _GEN_981; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire  _GEN_991 = deq_idxs_0[5] ? ~hit_tail_mask_0 : _GEN_984; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 105:44]
  wire [3:0] _GEN_992 = deq_idxs_0[5] ? fetch_buffer_5_gh_backup : _GEN_985; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire [31:0] _GEN_993 = deq_idxs_0[5] ? fetch_buffer_5_inst_addr : _GEN_986; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire [31:0] _GEN_994 = deq_idxs_0[5] ? fetch_buffer_5_inst : _GEN_987; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire  _GEN_995 = deq_idxs_0[6] ? fetch_buffer_6_predict_taken : _GEN_988; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire  _GEN_998 = deq_idxs_0[6] ? ~hit_tail_mask_0 : _GEN_991; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 105:44]
  wire [3:0] _GEN_999 = deq_idxs_0[6] ? fetch_buffer_6_gh_backup : _GEN_992; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire [31:0] _GEN_1000 = deq_idxs_0[6] ? fetch_buffer_6_inst_addr : _GEN_993; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire [31:0] _GEN_1001 = deq_idxs_0[6] ? fetch_buffer_6_inst : _GEN_994; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire  _GEN_1002 = deq_idxs_0[7] ? fetch_buffer_7_predict_taken : _GEN_995; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire  _GEN_1005 = deq_idxs_0[7] ? ~hit_tail_mask_0 : _GEN_998; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 105:44]
  wire [3:0] _GEN_1006 = deq_idxs_0[7] ? fetch_buffer_7_gh_backup : _GEN_999; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire [31:0] _GEN_1007 = deq_idxs_0[7] ? fetch_buffer_7_inst_addr : _GEN_1000; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire [31:0] _GEN_1008 = deq_idxs_0[7] ? fetch_buffer_7_inst : _GEN_1001; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire  _GEN_1009 = deq_idxs_0[8] ? fetch_buffer_8_predict_taken : _GEN_1002; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire  _GEN_1012 = deq_idxs_0[8] ? ~hit_tail_mask_0 : _GEN_1005; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 105:44]
  wire [3:0] _GEN_1013 = deq_idxs_0[8] ? fetch_buffer_8_gh_backup : _GEN_1006; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire [31:0] _GEN_1014 = deq_idxs_0[8] ? fetch_buffer_8_inst_addr : _GEN_1007; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire [31:0] _GEN_1015 = deq_idxs_0[8] ? fetch_buffer_8_inst : _GEN_1008; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire  _GEN_1016 = deq_idxs_0[9] ? fetch_buffer_9_predict_taken : _GEN_1009; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire  _GEN_1019 = deq_idxs_0[9] ? ~hit_tail_mask_0 : _GEN_1012; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 105:44]
  wire [3:0] _GEN_1020 = deq_idxs_0[9] ? fetch_buffer_9_gh_backup : _GEN_1013; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire [31:0] _GEN_1021 = deq_idxs_0[9] ? fetch_buffer_9_inst_addr : _GEN_1014; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire [31:0] _GEN_1022 = deq_idxs_0[9] ? fetch_buffer_9_inst : _GEN_1015; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire  _GEN_1023 = deq_idxs_0[10] ? fetch_buffer_10_predict_taken : _GEN_1016; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire  _GEN_1026 = deq_idxs_0[10] ? ~hit_tail_mask_0 : _GEN_1019; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 105:44]
  wire [3:0] _GEN_1027 = deq_idxs_0[10] ? fetch_buffer_10_gh_backup : _GEN_1020; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire [31:0] _GEN_1028 = deq_idxs_0[10] ? fetch_buffer_10_inst_addr : _GEN_1021; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire [31:0] _GEN_1029 = deq_idxs_0[10] ? fetch_buffer_10_inst : _GEN_1022; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire  _GEN_1030 = deq_idxs_0[11] ? fetch_buffer_11_predict_taken : _GEN_1023; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire  _GEN_1033 = deq_idxs_0[11] ? ~hit_tail_mask_0 : _GEN_1026; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 105:44]
  wire [3:0] _GEN_1034 = deq_idxs_0[11] ? fetch_buffer_11_gh_backup : _GEN_1027; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire [31:0] _GEN_1035 = deq_idxs_0[11] ? fetch_buffer_11_inst_addr : _GEN_1028; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire [31:0] _GEN_1036 = deq_idxs_0[11] ? fetch_buffer_11_inst : _GEN_1029; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire  _GEN_1037 = deq_idxs_0[12] ? fetch_buffer_12_predict_taken : _GEN_1030; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire  _GEN_1040 = deq_idxs_0[12] ? ~hit_tail_mask_0 : _GEN_1033; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 105:44]
  wire [3:0] _GEN_1041 = deq_idxs_0[12] ? fetch_buffer_12_gh_backup : _GEN_1034; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire [31:0] _GEN_1042 = deq_idxs_0[12] ? fetch_buffer_12_inst_addr : _GEN_1035; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire [31:0] _GEN_1043 = deq_idxs_0[12] ? fetch_buffer_12_inst : _GEN_1036; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire  _GEN_1044 = deq_idxs_0[13] ? fetch_buffer_13_predict_taken : _GEN_1037; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire  _GEN_1047 = deq_idxs_0[13] ? ~hit_tail_mask_0 : _GEN_1040; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 105:44]
  wire [3:0] _GEN_1048 = deq_idxs_0[13] ? fetch_buffer_13_gh_backup : _GEN_1041; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire [31:0] _GEN_1049 = deq_idxs_0[13] ? fetch_buffer_13_inst_addr : _GEN_1042; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire [31:0] _GEN_1050 = deq_idxs_0[13] ? fetch_buffer_13_inst : _GEN_1043; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire  _GEN_1051 = deq_idxs_0[14] ? fetch_buffer_14_predict_taken : _GEN_1044; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire  _GEN_1054 = deq_idxs_0[14] ? ~hit_tail_mask_0 : _GEN_1047; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 105:44]
  wire [3:0] _GEN_1055 = deq_idxs_0[14] ? fetch_buffer_14_gh_backup : _GEN_1048; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire [31:0] _GEN_1056 = deq_idxs_0[14] ? fetch_buffer_14_inst_addr : _GEN_1049; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire [31:0] _GEN_1057 = deq_idxs_0[14] ? fetch_buffer_14_inst : _GEN_1050; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire  _GEN_1058 = deq_idxs_0[15] ? fetch_buffer_15_predict_taken : _GEN_1051; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire  _GEN_1061 = deq_idxs_0[15] ? ~hit_tail_mask_0 : _GEN_1054; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 105:44]
  wire [3:0] _GEN_1062 = deq_idxs_0[15] ? fetch_buffer_15_gh_backup : _GEN_1055; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire [31:0] _GEN_1063 = deq_idxs_0[15] ? fetch_buffer_15_inst_addr : _GEN_1056; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire [31:0] _GEN_1064 = deq_idxs_0[15] ? fetch_buffer_15_inst : _GEN_1057; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire  _GEN_1079 = deq_idxs_1[1] ? fetch_buffer_1_predict_taken : fetch_buffer_0_predict_taken; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire  _GEN_1082 = deq_idxs_1[1] ? ~deq_invalid_1 : ~deq_invalid_1; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 105:44]
  wire [3:0] _GEN_1083 = deq_idxs_1[1] ? fetch_buffer_1_gh_backup : fetch_buffer_0_gh_backup; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire [31:0] _GEN_1084 = deq_idxs_1[1] ? fetch_buffer_1_inst_addr : fetch_buffer_0_inst_addr; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire [31:0] _GEN_1085 = deq_idxs_1[1] ? fetch_buffer_1_inst : fetch_buffer_0_inst; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire  _GEN_1086 = deq_idxs_1[2] ? fetch_buffer_2_predict_taken : _GEN_1079; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire  _GEN_1089 = deq_idxs_1[2] ? ~deq_invalid_1 : _GEN_1082; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 105:44]
  wire [3:0] _GEN_1090 = deq_idxs_1[2] ? fetch_buffer_2_gh_backup : _GEN_1083; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire [31:0] _GEN_1091 = deq_idxs_1[2] ? fetch_buffer_2_inst_addr : _GEN_1084; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire [31:0] _GEN_1092 = deq_idxs_1[2] ? fetch_buffer_2_inst : _GEN_1085; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire  _GEN_1093 = deq_idxs_1[3] ? fetch_buffer_3_predict_taken : _GEN_1086; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire  _GEN_1096 = deq_idxs_1[3] ? ~deq_invalid_1 : _GEN_1089; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 105:44]
  wire [3:0] _GEN_1097 = deq_idxs_1[3] ? fetch_buffer_3_gh_backup : _GEN_1090; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire [31:0] _GEN_1098 = deq_idxs_1[3] ? fetch_buffer_3_inst_addr : _GEN_1091; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire [31:0] _GEN_1099 = deq_idxs_1[3] ? fetch_buffer_3_inst : _GEN_1092; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire  _GEN_1100 = deq_idxs_1[4] ? fetch_buffer_4_predict_taken : _GEN_1093; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire  _GEN_1103 = deq_idxs_1[4] ? ~deq_invalid_1 : _GEN_1096; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 105:44]
  wire [3:0] _GEN_1104 = deq_idxs_1[4] ? fetch_buffer_4_gh_backup : _GEN_1097; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire [31:0] _GEN_1105 = deq_idxs_1[4] ? fetch_buffer_4_inst_addr : _GEN_1098; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire [31:0] _GEN_1106 = deq_idxs_1[4] ? fetch_buffer_4_inst : _GEN_1099; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire  _GEN_1107 = deq_idxs_1[5] ? fetch_buffer_5_predict_taken : _GEN_1100; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire  _GEN_1110 = deq_idxs_1[5] ? ~deq_invalid_1 : _GEN_1103; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 105:44]
  wire [3:0] _GEN_1111 = deq_idxs_1[5] ? fetch_buffer_5_gh_backup : _GEN_1104; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire [31:0] _GEN_1112 = deq_idxs_1[5] ? fetch_buffer_5_inst_addr : _GEN_1105; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire [31:0] _GEN_1113 = deq_idxs_1[5] ? fetch_buffer_5_inst : _GEN_1106; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire  _GEN_1114 = deq_idxs_1[6] ? fetch_buffer_6_predict_taken : _GEN_1107; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire  _GEN_1117 = deq_idxs_1[6] ? ~deq_invalid_1 : _GEN_1110; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 105:44]
  wire [3:0] _GEN_1118 = deq_idxs_1[6] ? fetch_buffer_6_gh_backup : _GEN_1111; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire [31:0] _GEN_1119 = deq_idxs_1[6] ? fetch_buffer_6_inst_addr : _GEN_1112; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire [31:0] _GEN_1120 = deq_idxs_1[6] ? fetch_buffer_6_inst : _GEN_1113; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire  _GEN_1121 = deq_idxs_1[7] ? fetch_buffer_7_predict_taken : _GEN_1114; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire  _GEN_1124 = deq_idxs_1[7] ? ~deq_invalid_1 : _GEN_1117; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 105:44]
  wire [3:0] _GEN_1125 = deq_idxs_1[7] ? fetch_buffer_7_gh_backup : _GEN_1118; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire [31:0] _GEN_1126 = deq_idxs_1[7] ? fetch_buffer_7_inst_addr : _GEN_1119; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire [31:0] _GEN_1127 = deq_idxs_1[7] ? fetch_buffer_7_inst : _GEN_1120; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire  _GEN_1128 = deq_idxs_1[8] ? fetch_buffer_8_predict_taken : _GEN_1121; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire  _GEN_1131 = deq_idxs_1[8] ? ~deq_invalid_1 : _GEN_1124; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 105:44]
  wire [3:0] _GEN_1132 = deq_idxs_1[8] ? fetch_buffer_8_gh_backup : _GEN_1125; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire [31:0] _GEN_1133 = deq_idxs_1[8] ? fetch_buffer_8_inst_addr : _GEN_1126; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire [31:0] _GEN_1134 = deq_idxs_1[8] ? fetch_buffer_8_inst : _GEN_1127; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire  _GEN_1135 = deq_idxs_1[9] ? fetch_buffer_9_predict_taken : _GEN_1128; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire  _GEN_1138 = deq_idxs_1[9] ? ~deq_invalid_1 : _GEN_1131; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 105:44]
  wire [3:0] _GEN_1139 = deq_idxs_1[9] ? fetch_buffer_9_gh_backup : _GEN_1132; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire [31:0] _GEN_1140 = deq_idxs_1[9] ? fetch_buffer_9_inst_addr : _GEN_1133; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire [31:0] _GEN_1141 = deq_idxs_1[9] ? fetch_buffer_9_inst : _GEN_1134; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire  _GEN_1142 = deq_idxs_1[10] ? fetch_buffer_10_predict_taken : _GEN_1135; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire  _GEN_1145 = deq_idxs_1[10] ? ~deq_invalid_1 : _GEN_1138; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 105:44]
  wire [3:0] _GEN_1146 = deq_idxs_1[10] ? fetch_buffer_10_gh_backup : _GEN_1139; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire [31:0] _GEN_1147 = deq_idxs_1[10] ? fetch_buffer_10_inst_addr : _GEN_1140; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire [31:0] _GEN_1148 = deq_idxs_1[10] ? fetch_buffer_10_inst : _GEN_1141; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire  _GEN_1149 = deq_idxs_1[11] ? fetch_buffer_11_predict_taken : _GEN_1142; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire  _GEN_1152 = deq_idxs_1[11] ? ~deq_invalid_1 : _GEN_1145; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 105:44]
  wire [3:0] _GEN_1153 = deq_idxs_1[11] ? fetch_buffer_11_gh_backup : _GEN_1146; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire [31:0] _GEN_1154 = deq_idxs_1[11] ? fetch_buffer_11_inst_addr : _GEN_1147; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire [31:0] _GEN_1155 = deq_idxs_1[11] ? fetch_buffer_11_inst : _GEN_1148; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire  _GEN_1156 = deq_idxs_1[12] ? fetch_buffer_12_predict_taken : _GEN_1149; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire  _GEN_1159 = deq_idxs_1[12] ? ~deq_invalid_1 : _GEN_1152; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 105:44]
  wire [3:0] _GEN_1160 = deq_idxs_1[12] ? fetch_buffer_12_gh_backup : _GEN_1153; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire [31:0] _GEN_1161 = deq_idxs_1[12] ? fetch_buffer_12_inst_addr : _GEN_1154; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire [31:0] _GEN_1162 = deq_idxs_1[12] ? fetch_buffer_12_inst : _GEN_1155; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire  _GEN_1163 = deq_idxs_1[13] ? fetch_buffer_13_predict_taken : _GEN_1156; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire  _GEN_1166 = deq_idxs_1[13] ? ~deq_invalid_1 : _GEN_1159; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 105:44]
  wire [3:0] _GEN_1167 = deq_idxs_1[13] ? fetch_buffer_13_gh_backup : _GEN_1160; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire [31:0] _GEN_1168 = deq_idxs_1[13] ? fetch_buffer_13_inst_addr : _GEN_1161; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire [31:0] _GEN_1169 = deq_idxs_1[13] ? fetch_buffer_13_inst : _GEN_1162; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire  _GEN_1170 = deq_idxs_1[14] ? fetch_buffer_14_predict_taken : _GEN_1163; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire  _GEN_1173 = deq_idxs_1[14] ? ~deq_invalid_1 : _GEN_1166; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 105:44]
  wire [3:0] _GEN_1174 = deq_idxs_1[14] ? fetch_buffer_14_gh_backup : _GEN_1167; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire [31:0] _GEN_1175 = deq_idxs_1[14] ? fetch_buffer_14_inst_addr : _GEN_1168; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire [31:0] _GEN_1176 = deq_idxs_1[14] ? fetch_buffer_14_inst : _GEN_1169; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire  _GEN_1177 = deq_idxs_1[15] ? fetch_buffer_15_predict_taken : _GEN_1170; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire  _GEN_1180 = deq_idxs_1[15] ? ~deq_invalid_1 : _GEN_1173; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 105:44]
  wire [3:0] _GEN_1181 = deq_idxs_1[15] ? fetch_buffer_15_gh_backup : _GEN_1174; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire [31:0] _GEN_1182 = deq_idxs_1[15] ? fetch_buffer_15_inst_addr : _GEN_1175; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire [31:0] _GEN_1183 = deq_idxs_1[15] ? fetch_buffer_15_inst : _GEN_1176; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  wire [16:0] _T_458 = io_fb_resp_deq_valid_0 ? deq_idxs_1 : deq_idxs_0; // @[FetchBuffer.scala 111:20]
  wire [15:0] hi_9 = _T_458[15:0]; // @[FetchBuffer.scala 42:12]
  wire  lo_9 = _T_458[16]; // @[FetchBuffer.scala 42:29]
  wire [16:0] _T_459 = {hi_9,lo_9}; // @[Cat.scala 30:58]
  wire  _GEN_1191 = do_enq | maybe_full; // @[FetchBuffer.scala 121:22 FetchBuffer.scala 122:16 FetchBuffer.scala 53:29]
  wire  _GEN_1192 = do_deq ? 1'h0 : _GEN_1191; // @[FetchBuffer.scala 119:22 FetchBuffer.scala 120:16]
  wire  _GEN_1193 = do_deq & do_enq | _GEN_1192; // @[FetchBuffer.scala 117:26 FetchBuffer.scala 118:16]
  assign io_bpu_inst_packet_i_ready = _do_enq_T_2 | ~io_bpu_inst_packet_i_valid | ~_do_enq_T_10; // @[FetchBuffer.scala 131:105]
  assign io_inst_bank_valid = ~is_empty & ~io_clear_i; // @[FetchBuffer.scala 115:35]
  assign io_inst_bank_bits_data_0_inst = deq_idxs_lo ? fetch_buffer_16_inst : _GEN_1064; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  assign io_inst_bank_bits_data_0_inst_addr = deq_idxs_lo ? fetch_buffer_16_inst_addr : _GEN_1063; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  assign io_inst_bank_bits_data_0_gh_backup = deq_idxs_lo ? fetch_buffer_16_gh_backup : _GEN_1062; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  assign io_inst_bank_bits_data_0_is_valid = deq_idxs_lo ? ~hit_tail_mask_0 : _GEN_1061; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 105:44]
  assign io_inst_bank_bits_data_0_predict_taken = deq_idxs_lo ? fetch_buffer_16_predict_taken : _GEN_1058; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  assign io_inst_bank_bits_data_1_inst = deq_idxs_1[16] ? fetch_buffer_16_inst : _GEN_1183; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  assign io_inst_bank_bits_data_1_inst_addr = deq_idxs_1[16] ? fetch_buffer_16_inst_addr : _GEN_1182; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  assign io_inst_bank_bits_data_1_gh_backup = deq_idxs_1[16] ? fetch_buffer_16_gh_backup : _GEN_1181; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  assign io_inst_bank_bits_data_1_is_valid = deq_idxs_1[16] ? ~deq_invalid_1 : _GEN_1180; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 105:44]
  assign io_inst_bank_bits_data_1_predict_taken = deq_idxs_1[16] ? fetch_buffer_16_predict_taken : _GEN_1177; // @[FetchBuffer.scala 103:28 FetchBuffer.scala 104:35]
  always @(posedge clock) begin
    if (reset) begin // @[FetchBuffer.scala 134:24]
      fetch_buffer_0_inst <= 32'h0; // @[FetchBuffer.scala 17:19]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_7 & enq_idxs_7[0]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_0_inst <= io_bpu_inst_packet_i_bits_data_7; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_6 & enq_idxs_6[0]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_0_inst <= io_bpu_inst_packet_i_bits_data_6; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_5 & enq_idxs_5[0]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_0_inst <= io_bpu_inst_packet_i_bits_data_5; // @[FetchBuffer.scala 85:25]
    end else begin
      fetch_buffer_0_inst <= _GEN_482;
    end
    if (reset) begin // @[FetchBuffer.scala 134:24]
      fetch_buffer_0_inst_addr <= 32'h0; // @[FetchBuffer.scala 18:19]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_7 & enq_idxs_7[0]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_0_inst_addr <= inst_packet_7_inst_addr; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_6 & enq_idxs_6[0]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_0_inst_addr <= inst_packet_6_inst_addr; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_5 & enq_idxs_5[0]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_0_inst_addr <= inst_packet_5_inst_addr; // @[FetchBuffer.scala 85:25]
    end else begin
      fetch_buffer_0_inst_addr <= _GEN_481;
    end
    if (reset) begin // @[FetchBuffer.scala 134:24]
      fetch_buffer_0_gh_backup <= 4'h0; // @[FetchBuffer.scala 19:19]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_7 & enq_idxs_7[0]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_0_gh_backup <= io_bpu_inst_packet_i_bits_gh_backup; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_6 & enq_idxs_6[0]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_0_gh_backup <= io_bpu_inst_packet_i_bits_gh_backup; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_5 & enq_idxs_5[0]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_0_gh_backup <= io_bpu_inst_packet_i_bits_gh_backup; // @[FetchBuffer.scala 85:25]
    end else begin
      fetch_buffer_0_gh_backup <= _GEN_480;
    end
    if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_7 & enq_idxs_7[0]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_0_predict_taken <= io_bpu_inst_packet_i_bits_predict_mask_7; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_6 & enq_idxs_6[0]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_0_predict_taken <= io_bpu_inst_packet_i_bits_predict_mask_6; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_5 & enq_idxs_5[0]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_0_predict_taken <= io_bpu_inst_packet_i_bits_predict_mask_5; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_4 & enq_idxs_4[0]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_0_predict_taken <= io_bpu_inst_packet_i_bits_predict_mask_4; // @[FetchBuffer.scala 85:25]
    end else begin
      fetch_buffer_0_predict_taken <= _GEN_357;
    end
    if (reset) begin // @[FetchBuffer.scala 134:24]
      fetch_buffer_1_inst <= 32'h0; // @[FetchBuffer.scala 17:19]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_7 & enq_idxs_7[1]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_1_inst <= io_bpu_inst_packet_i_bits_data_7; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_6 & enq_idxs_6[1]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_1_inst <= io_bpu_inst_packet_i_bits_data_6; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_5 & enq_idxs_5[1]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_1_inst <= io_bpu_inst_packet_i_bits_data_5; // @[FetchBuffer.scala 85:25]
    end else begin
      fetch_buffer_1_inst <= _GEN_489;
    end
    if (reset) begin // @[FetchBuffer.scala 134:24]
      fetch_buffer_1_inst_addr <= 32'h0; // @[FetchBuffer.scala 18:19]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_7 & enq_idxs_7[1]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_1_inst_addr <= inst_packet_7_inst_addr; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_6 & enq_idxs_6[1]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_1_inst_addr <= inst_packet_6_inst_addr; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_5 & enq_idxs_5[1]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_1_inst_addr <= inst_packet_5_inst_addr; // @[FetchBuffer.scala 85:25]
    end else begin
      fetch_buffer_1_inst_addr <= _GEN_488;
    end
    if (reset) begin // @[FetchBuffer.scala 134:24]
      fetch_buffer_1_gh_backup <= 4'h0; // @[FetchBuffer.scala 19:19]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_7 & enq_idxs_7[1]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_1_gh_backup <= io_bpu_inst_packet_i_bits_gh_backup; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_6 & enq_idxs_6[1]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_1_gh_backup <= io_bpu_inst_packet_i_bits_gh_backup; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_5 & enq_idxs_5[1]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_1_gh_backup <= io_bpu_inst_packet_i_bits_gh_backup; // @[FetchBuffer.scala 85:25]
    end else begin
      fetch_buffer_1_gh_backup <= _GEN_487;
    end
    if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_7 & enq_idxs_7[1]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_1_predict_taken <= io_bpu_inst_packet_i_bits_predict_mask_7; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_6 & enq_idxs_6[1]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_1_predict_taken <= io_bpu_inst_packet_i_bits_predict_mask_6; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_5 & enq_idxs_5[1]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_1_predict_taken <= io_bpu_inst_packet_i_bits_predict_mask_5; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_4 & enq_idxs_4[1]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_1_predict_taken <= io_bpu_inst_packet_i_bits_predict_mask_4; // @[FetchBuffer.scala 85:25]
    end else begin
      fetch_buffer_1_predict_taken <= _GEN_364;
    end
    if (reset) begin // @[FetchBuffer.scala 134:24]
      fetch_buffer_2_inst <= 32'h0; // @[FetchBuffer.scala 17:19]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_7 & enq_idxs_7[2]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_2_inst <= io_bpu_inst_packet_i_bits_data_7; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_6 & enq_idxs_6[2]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_2_inst <= io_bpu_inst_packet_i_bits_data_6; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_5 & enq_idxs_5[2]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_2_inst <= io_bpu_inst_packet_i_bits_data_5; // @[FetchBuffer.scala 85:25]
    end else begin
      fetch_buffer_2_inst <= _GEN_496;
    end
    if (reset) begin // @[FetchBuffer.scala 134:24]
      fetch_buffer_2_inst_addr <= 32'h0; // @[FetchBuffer.scala 18:19]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_7 & enq_idxs_7[2]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_2_inst_addr <= inst_packet_7_inst_addr; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_6 & enq_idxs_6[2]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_2_inst_addr <= inst_packet_6_inst_addr; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_5 & enq_idxs_5[2]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_2_inst_addr <= inst_packet_5_inst_addr; // @[FetchBuffer.scala 85:25]
    end else begin
      fetch_buffer_2_inst_addr <= _GEN_495;
    end
    if (reset) begin // @[FetchBuffer.scala 134:24]
      fetch_buffer_2_gh_backup <= 4'h0; // @[FetchBuffer.scala 19:19]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_7 & enq_idxs_7[2]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_2_gh_backup <= io_bpu_inst_packet_i_bits_gh_backup; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_6 & enq_idxs_6[2]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_2_gh_backup <= io_bpu_inst_packet_i_bits_gh_backup; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_5 & enq_idxs_5[2]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_2_gh_backup <= io_bpu_inst_packet_i_bits_gh_backup; // @[FetchBuffer.scala 85:25]
    end else begin
      fetch_buffer_2_gh_backup <= _GEN_494;
    end
    if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_7 & enq_idxs_7[2]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_2_predict_taken <= io_bpu_inst_packet_i_bits_predict_mask_7; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_6 & enq_idxs_6[2]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_2_predict_taken <= io_bpu_inst_packet_i_bits_predict_mask_6; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_5 & enq_idxs_5[2]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_2_predict_taken <= io_bpu_inst_packet_i_bits_predict_mask_5; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_4 & enq_idxs_4[2]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_2_predict_taken <= io_bpu_inst_packet_i_bits_predict_mask_4; // @[FetchBuffer.scala 85:25]
    end else begin
      fetch_buffer_2_predict_taken <= _GEN_371;
    end
    if (reset) begin // @[FetchBuffer.scala 134:24]
      fetch_buffer_3_inst <= 32'h0; // @[FetchBuffer.scala 17:19]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_7 & enq_idxs_7[3]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_3_inst <= io_bpu_inst_packet_i_bits_data_7; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_6 & enq_idxs_6[3]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_3_inst <= io_bpu_inst_packet_i_bits_data_6; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_5 & enq_idxs_5[3]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_3_inst <= io_bpu_inst_packet_i_bits_data_5; // @[FetchBuffer.scala 85:25]
    end else begin
      fetch_buffer_3_inst <= _GEN_503;
    end
    if (reset) begin // @[FetchBuffer.scala 134:24]
      fetch_buffer_3_inst_addr <= 32'h0; // @[FetchBuffer.scala 18:19]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_7 & enq_idxs_7[3]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_3_inst_addr <= inst_packet_7_inst_addr; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_6 & enq_idxs_6[3]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_3_inst_addr <= inst_packet_6_inst_addr; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_5 & enq_idxs_5[3]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_3_inst_addr <= inst_packet_5_inst_addr; // @[FetchBuffer.scala 85:25]
    end else begin
      fetch_buffer_3_inst_addr <= _GEN_502;
    end
    if (reset) begin // @[FetchBuffer.scala 134:24]
      fetch_buffer_3_gh_backup <= 4'h0; // @[FetchBuffer.scala 19:19]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_7 & enq_idxs_7[3]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_3_gh_backup <= io_bpu_inst_packet_i_bits_gh_backup; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_6 & enq_idxs_6[3]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_3_gh_backup <= io_bpu_inst_packet_i_bits_gh_backup; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_5 & enq_idxs_5[3]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_3_gh_backup <= io_bpu_inst_packet_i_bits_gh_backup; // @[FetchBuffer.scala 85:25]
    end else begin
      fetch_buffer_3_gh_backup <= _GEN_501;
    end
    if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_7 & enq_idxs_7[3]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_3_predict_taken <= io_bpu_inst_packet_i_bits_predict_mask_7; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_6 & enq_idxs_6[3]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_3_predict_taken <= io_bpu_inst_packet_i_bits_predict_mask_6; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_5 & enq_idxs_5[3]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_3_predict_taken <= io_bpu_inst_packet_i_bits_predict_mask_5; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_4 & enq_idxs_4[3]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_3_predict_taken <= io_bpu_inst_packet_i_bits_predict_mask_4; // @[FetchBuffer.scala 85:25]
    end else begin
      fetch_buffer_3_predict_taken <= _GEN_378;
    end
    if (reset) begin // @[FetchBuffer.scala 134:24]
      fetch_buffer_4_inst <= 32'h0; // @[FetchBuffer.scala 17:19]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_7 & enq_idxs_7[4]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_4_inst <= io_bpu_inst_packet_i_bits_data_7; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_6 & enq_idxs_6[4]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_4_inst <= io_bpu_inst_packet_i_bits_data_6; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_5 & enq_idxs_5[4]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_4_inst <= io_bpu_inst_packet_i_bits_data_5; // @[FetchBuffer.scala 85:25]
    end else begin
      fetch_buffer_4_inst <= _GEN_510;
    end
    if (reset) begin // @[FetchBuffer.scala 134:24]
      fetch_buffer_4_inst_addr <= 32'h0; // @[FetchBuffer.scala 18:19]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_7 & enq_idxs_7[4]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_4_inst_addr <= inst_packet_7_inst_addr; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_6 & enq_idxs_6[4]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_4_inst_addr <= inst_packet_6_inst_addr; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_5 & enq_idxs_5[4]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_4_inst_addr <= inst_packet_5_inst_addr; // @[FetchBuffer.scala 85:25]
    end else begin
      fetch_buffer_4_inst_addr <= _GEN_509;
    end
    if (reset) begin // @[FetchBuffer.scala 134:24]
      fetch_buffer_4_gh_backup <= 4'h0; // @[FetchBuffer.scala 19:19]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_7 & enq_idxs_7[4]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_4_gh_backup <= io_bpu_inst_packet_i_bits_gh_backup; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_6 & enq_idxs_6[4]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_4_gh_backup <= io_bpu_inst_packet_i_bits_gh_backup; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_5 & enq_idxs_5[4]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_4_gh_backup <= io_bpu_inst_packet_i_bits_gh_backup; // @[FetchBuffer.scala 85:25]
    end else begin
      fetch_buffer_4_gh_backup <= _GEN_508;
    end
    if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_7 & enq_idxs_7[4]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_4_predict_taken <= io_bpu_inst_packet_i_bits_predict_mask_7; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_6 & enq_idxs_6[4]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_4_predict_taken <= io_bpu_inst_packet_i_bits_predict_mask_6; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_5 & enq_idxs_5[4]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_4_predict_taken <= io_bpu_inst_packet_i_bits_predict_mask_5; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_4 & enq_idxs_4[4]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_4_predict_taken <= io_bpu_inst_packet_i_bits_predict_mask_4; // @[FetchBuffer.scala 85:25]
    end else begin
      fetch_buffer_4_predict_taken <= _GEN_385;
    end
    if (reset) begin // @[FetchBuffer.scala 134:24]
      fetch_buffer_5_inst <= 32'h0; // @[FetchBuffer.scala 17:19]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_7 & enq_idxs_7[5]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_5_inst <= io_bpu_inst_packet_i_bits_data_7; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_6 & enq_idxs_6[5]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_5_inst <= io_bpu_inst_packet_i_bits_data_6; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_5 & enq_idxs_5[5]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_5_inst <= io_bpu_inst_packet_i_bits_data_5; // @[FetchBuffer.scala 85:25]
    end else begin
      fetch_buffer_5_inst <= _GEN_517;
    end
    if (reset) begin // @[FetchBuffer.scala 134:24]
      fetch_buffer_5_inst_addr <= 32'h0; // @[FetchBuffer.scala 18:19]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_7 & enq_idxs_7[5]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_5_inst_addr <= inst_packet_7_inst_addr; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_6 & enq_idxs_6[5]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_5_inst_addr <= inst_packet_6_inst_addr; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_5 & enq_idxs_5[5]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_5_inst_addr <= inst_packet_5_inst_addr; // @[FetchBuffer.scala 85:25]
    end else begin
      fetch_buffer_5_inst_addr <= _GEN_516;
    end
    if (reset) begin // @[FetchBuffer.scala 134:24]
      fetch_buffer_5_gh_backup <= 4'h0; // @[FetchBuffer.scala 19:19]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_7 & enq_idxs_7[5]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_5_gh_backup <= io_bpu_inst_packet_i_bits_gh_backup; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_6 & enq_idxs_6[5]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_5_gh_backup <= io_bpu_inst_packet_i_bits_gh_backup; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_5 & enq_idxs_5[5]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_5_gh_backup <= io_bpu_inst_packet_i_bits_gh_backup; // @[FetchBuffer.scala 85:25]
    end else begin
      fetch_buffer_5_gh_backup <= _GEN_515;
    end
    if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_7 & enq_idxs_7[5]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_5_predict_taken <= io_bpu_inst_packet_i_bits_predict_mask_7; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_6 & enq_idxs_6[5]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_5_predict_taken <= io_bpu_inst_packet_i_bits_predict_mask_6; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_5 & enq_idxs_5[5]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_5_predict_taken <= io_bpu_inst_packet_i_bits_predict_mask_5; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_4 & enq_idxs_4[5]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_5_predict_taken <= io_bpu_inst_packet_i_bits_predict_mask_4; // @[FetchBuffer.scala 85:25]
    end else begin
      fetch_buffer_5_predict_taken <= _GEN_392;
    end
    if (reset) begin // @[FetchBuffer.scala 134:24]
      fetch_buffer_6_inst <= 32'h0; // @[FetchBuffer.scala 17:19]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_7 & enq_idxs_7[6]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_6_inst <= io_bpu_inst_packet_i_bits_data_7; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_6 & enq_idxs_6[6]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_6_inst <= io_bpu_inst_packet_i_bits_data_6; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_5 & enq_idxs_5[6]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_6_inst <= io_bpu_inst_packet_i_bits_data_5; // @[FetchBuffer.scala 85:25]
    end else begin
      fetch_buffer_6_inst <= _GEN_524;
    end
    if (reset) begin // @[FetchBuffer.scala 134:24]
      fetch_buffer_6_inst_addr <= 32'h0; // @[FetchBuffer.scala 18:19]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_7 & enq_idxs_7[6]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_6_inst_addr <= inst_packet_7_inst_addr; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_6 & enq_idxs_6[6]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_6_inst_addr <= inst_packet_6_inst_addr; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_5 & enq_idxs_5[6]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_6_inst_addr <= inst_packet_5_inst_addr; // @[FetchBuffer.scala 85:25]
    end else begin
      fetch_buffer_6_inst_addr <= _GEN_523;
    end
    if (reset) begin // @[FetchBuffer.scala 134:24]
      fetch_buffer_6_gh_backup <= 4'h0; // @[FetchBuffer.scala 19:19]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_7 & enq_idxs_7[6]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_6_gh_backup <= io_bpu_inst_packet_i_bits_gh_backup; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_6 & enq_idxs_6[6]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_6_gh_backup <= io_bpu_inst_packet_i_bits_gh_backup; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_5 & enq_idxs_5[6]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_6_gh_backup <= io_bpu_inst_packet_i_bits_gh_backup; // @[FetchBuffer.scala 85:25]
    end else begin
      fetch_buffer_6_gh_backup <= _GEN_522;
    end
    if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_7 & enq_idxs_7[6]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_6_predict_taken <= io_bpu_inst_packet_i_bits_predict_mask_7; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_6 & enq_idxs_6[6]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_6_predict_taken <= io_bpu_inst_packet_i_bits_predict_mask_6; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_5 & enq_idxs_5[6]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_6_predict_taken <= io_bpu_inst_packet_i_bits_predict_mask_5; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_4 & enq_idxs_4[6]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_6_predict_taken <= io_bpu_inst_packet_i_bits_predict_mask_4; // @[FetchBuffer.scala 85:25]
    end else begin
      fetch_buffer_6_predict_taken <= _GEN_399;
    end
    if (reset) begin // @[FetchBuffer.scala 134:24]
      fetch_buffer_7_inst <= 32'h0; // @[FetchBuffer.scala 17:19]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_7 & enq_idxs_7[7]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_7_inst <= io_bpu_inst_packet_i_bits_data_7; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_6 & enq_idxs_6[7]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_7_inst <= io_bpu_inst_packet_i_bits_data_6; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_5 & enq_idxs_5[7]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_7_inst <= io_bpu_inst_packet_i_bits_data_5; // @[FetchBuffer.scala 85:25]
    end else begin
      fetch_buffer_7_inst <= _GEN_531;
    end
    if (reset) begin // @[FetchBuffer.scala 134:24]
      fetch_buffer_7_inst_addr <= 32'h0; // @[FetchBuffer.scala 18:19]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_7 & enq_idxs_7[7]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_7_inst_addr <= inst_packet_7_inst_addr; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_6 & enq_idxs_6[7]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_7_inst_addr <= inst_packet_6_inst_addr; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_5 & enq_idxs_5[7]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_7_inst_addr <= inst_packet_5_inst_addr; // @[FetchBuffer.scala 85:25]
    end else begin
      fetch_buffer_7_inst_addr <= _GEN_530;
    end
    if (reset) begin // @[FetchBuffer.scala 134:24]
      fetch_buffer_7_gh_backup <= 4'h0; // @[FetchBuffer.scala 19:19]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_7 & enq_idxs_7[7]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_7_gh_backup <= io_bpu_inst_packet_i_bits_gh_backup; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_6 & enq_idxs_6[7]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_7_gh_backup <= io_bpu_inst_packet_i_bits_gh_backup; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_5 & enq_idxs_5[7]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_7_gh_backup <= io_bpu_inst_packet_i_bits_gh_backup; // @[FetchBuffer.scala 85:25]
    end else begin
      fetch_buffer_7_gh_backup <= _GEN_529;
    end
    if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_7 & enq_idxs_7[7]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_7_predict_taken <= io_bpu_inst_packet_i_bits_predict_mask_7; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_6 & enq_idxs_6[7]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_7_predict_taken <= io_bpu_inst_packet_i_bits_predict_mask_6; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_5 & enq_idxs_5[7]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_7_predict_taken <= io_bpu_inst_packet_i_bits_predict_mask_5; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_4 & enq_idxs_4[7]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_7_predict_taken <= io_bpu_inst_packet_i_bits_predict_mask_4; // @[FetchBuffer.scala 85:25]
    end else begin
      fetch_buffer_7_predict_taken <= _GEN_406;
    end
    if (reset) begin // @[FetchBuffer.scala 134:24]
      fetch_buffer_8_inst <= 32'h0; // @[FetchBuffer.scala 17:19]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_7 & enq_idxs_7[8]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_8_inst <= io_bpu_inst_packet_i_bits_data_7; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_6 & enq_idxs_6[8]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_8_inst <= io_bpu_inst_packet_i_bits_data_6; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_5 & enq_idxs_5[8]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_8_inst <= io_bpu_inst_packet_i_bits_data_5; // @[FetchBuffer.scala 85:25]
    end else begin
      fetch_buffer_8_inst <= _GEN_538;
    end
    if (reset) begin // @[FetchBuffer.scala 134:24]
      fetch_buffer_8_inst_addr <= 32'h0; // @[FetchBuffer.scala 18:19]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_7 & enq_idxs_7[8]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_8_inst_addr <= inst_packet_7_inst_addr; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_6 & enq_idxs_6[8]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_8_inst_addr <= inst_packet_6_inst_addr; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_5 & enq_idxs_5[8]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_8_inst_addr <= inst_packet_5_inst_addr; // @[FetchBuffer.scala 85:25]
    end else begin
      fetch_buffer_8_inst_addr <= _GEN_537;
    end
    if (reset) begin // @[FetchBuffer.scala 134:24]
      fetch_buffer_8_gh_backup <= 4'h0; // @[FetchBuffer.scala 19:19]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_7 & enq_idxs_7[8]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_8_gh_backup <= io_bpu_inst_packet_i_bits_gh_backup; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_6 & enq_idxs_6[8]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_8_gh_backup <= io_bpu_inst_packet_i_bits_gh_backup; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_5 & enq_idxs_5[8]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_8_gh_backup <= io_bpu_inst_packet_i_bits_gh_backup; // @[FetchBuffer.scala 85:25]
    end else begin
      fetch_buffer_8_gh_backup <= _GEN_536;
    end
    if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_7 & enq_idxs_7[8]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_8_predict_taken <= io_bpu_inst_packet_i_bits_predict_mask_7; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_6 & enq_idxs_6[8]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_8_predict_taken <= io_bpu_inst_packet_i_bits_predict_mask_6; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_5 & enq_idxs_5[8]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_8_predict_taken <= io_bpu_inst_packet_i_bits_predict_mask_5; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_4 & enq_idxs_4[8]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_8_predict_taken <= io_bpu_inst_packet_i_bits_predict_mask_4; // @[FetchBuffer.scala 85:25]
    end else begin
      fetch_buffer_8_predict_taken <= _GEN_413;
    end
    if (reset) begin // @[FetchBuffer.scala 134:24]
      fetch_buffer_9_inst <= 32'h0; // @[FetchBuffer.scala 17:19]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_7 & enq_idxs_7[9]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_9_inst <= io_bpu_inst_packet_i_bits_data_7; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_6 & enq_idxs_6[9]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_9_inst <= io_bpu_inst_packet_i_bits_data_6; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_5 & enq_idxs_5[9]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_9_inst <= io_bpu_inst_packet_i_bits_data_5; // @[FetchBuffer.scala 85:25]
    end else begin
      fetch_buffer_9_inst <= _GEN_545;
    end
    if (reset) begin // @[FetchBuffer.scala 134:24]
      fetch_buffer_9_inst_addr <= 32'h0; // @[FetchBuffer.scala 18:19]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_7 & enq_idxs_7[9]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_9_inst_addr <= inst_packet_7_inst_addr; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_6 & enq_idxs_6[9]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_9_inst_addr <= inst_packet_6_inst_addr; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_5 & enq_idxs_5[9]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_9_inst_addr <= inst_packet_5_inst_addr; // @[FetchBuffer.scala 85:25]
    end else begin
      fetch_buffer_9_inst_addr <= _GEN_544;
    end
    if (reset) begin // @[FetchBuffer.scala 134:24]
      fetch_buffer_9_gh_backup <= 4'h0; // @[FetchBuffer.scala 19:19]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_7 & enq_idxs_7[9]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_9_gh_backup <= io_bpu_inst_packet_i_bits_gh_backup; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_6 & enq_idxs_6[9]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_9_gh_backup <= io_bpu_inst_packet_i_bits_gh_backup; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_5 & enq_idxs_5[9]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_9_gh_backup <= io_bpu_inst_packet_i_bits_gh_backup; // @[FetchBuffer.scala 85:25]
    end else begin
      fetch_buffer_9_gh_backup <= _GEN_543;
    end
    if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_7 & enq_idxs_7[9]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_9_predict_taken <= io_bpu_inst_packet_i_bits_predict_mask_7; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_6 & enq_idxs_6[9]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_9_predict_taken <= io_bpu_inst_packet_i_bits_predict_mask_6; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_5 & enq_idxs_5[9]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_9_predict_taken <= io_bpu_inst_packet_i_bits_predict_mask_5; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_4 & enq_idxs_4[9]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_9_predict_taken <= io_bpu_inst_packet_i_bits_predict_mask_4; // @[FetchBuffer.scala 85:25]
    end else begin
      fetch_buffer_9_predict_taken <= _GEN_420;
    end
    if (reset) begin // @[FetchBuffer.scala 134:24]
      fetch_buffer_10_inst <= 32'h0; // @[FetchBuffer.scala 17:19]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_7 & enq_idxs_7[10]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_10_inst <= io_bpu_inst_packet_i_bits_data_7; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_6 & enq_idxs_6[10]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_10_inst <= io_bpu_inst_packet_i_bits_data_6; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_5 & enq_idxs_5[10]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_10_inst <= io_bpu_inst_packet_i_bits_data_5; // @[FetchBuffer.scala 85:25]
    end else begin
      fetch_buffer_10_inst <= _GEN_552;
    end
    if (reset) begin // @[FetchBuffer.scala 134:24]
      fetch_buffer_10_inst_addr <= 32'h0; // @[FetchBuffer.scala 18:19]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_7 & enq_idxs_7[10]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_10_inst_addr <= inst_packet_7_inst_addr; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_6 & enq_idxs_6[10]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_10_inst_addr <= inst_packet_6_inst_addr; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_5 & enq_idxs_5[10]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_10_inst_addr <= inst_packet_5_inst_addr; // @[FetchBuffer.scala 85:25]
    end else begin
      fetch_buffer_10_inst_addr <= _GEN_551;
    end
    if (reset) begin // @[FetchBuffer.scala 134:24]
      fetch_buffer_10_gh_backup <= 4'h0; // @[FetchBuffer.scala 19:19]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_7 & enq_idxs_7[10]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_10_gh_backup <= io_bpu_inst_packet_i_bits_gh_backup; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_6 & enq_idxs_6[10]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_10_gh_backup <= io_bpu_inst_packet_i_bits_gh_backup; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_5 & enq_idxs_5[10]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_10_gh_backup <= io_bpu_inst_packet_i_bits_gh_backup; // @[FetchBuffer.scala 85:25]
    end else begin
      fetch_buffer_10_gh_backup <= _GEN_550;
    end
    if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_7 & enq_idxs_7[10]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_10_predict_taken <= io_bpu_inst_packet_i_bits_predict_mask_7; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_6 & enq_idxs_6[10]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_10_predict_taken <= io_bpu_inst_packet_i_bits_predict_mask_6; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_5 & enq_idxs_5[10]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_10_predict_taken <= io_bpu_inst_packet_i_bits_predict_mask_5; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_4 & enq_idxs_4[10]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_10_predict_taken <= io_bpu_inst_packet_i_bits_predict_mask_4; // @[FetchBuffer.scala 85:25]
    end else begin
      fetch_buffer_10_predict_taken <= _GEN_427;
    end
    if (reset) begin // @[FetchBuffer.scala 134:24]
      fetch_buffer_11_inst <= 32'h0; // @[FetchBuffer.scala 17:19]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_7 & enq_idxs_7[11]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_11_inst <= io_bpu_inst_packet_i_bits_data_7; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_6 & enq_idxs_6[11]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_11_inst <= io_bpu_inst_packet_i_bits_data_6; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_5 & enq_idxs_5[11]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_11_inst <= io_bpu_inst_packet_i_bits_data_5; // @[FetchBuffer.scala 85:25]
    end else begin
      fetch_buffer_11_inst <= _GEN_559;
    end
    if (reset) begin // @[FetchBuffer.scala 134:24]
      fetch_buffer_11_inst_addr <= 32'h0; // @[FetchBuffer.scala 18:19]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_7 & enq_idxs_7[11]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_11_inst_addr <= inst_packet_7_inst_addr; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_6 & enq_idxs_6[11]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_11_inst_addr <= inst_packet_6_inst_addr; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_5 & enq_idxs_5[11]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_11_inst_addr <= inst_packet_5_inst_addr; // @[FetchBuffer.scala 85:25]
    end else begin
      fetch_buffer_11_inst_addr <= _GEN_558;
    end
    if (reset) begin // @[FetchBuffer.scala 134:24]
      fetch_buffer_11_gh_backup <= 4'h0; // @[FetchBuffer.scala 19:19]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_7 & enq_idxs_7[11]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_11_gh_backup <= io_bpu_inst_packet_i_bits_gh_backup; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_6 & enq_idxs_6[11]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_11_gh_backup <= io_bpu_inst_packet_i_bits_gh_backup; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_5 & enq_idxs_5[11]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_11_gh_backup <= io_bpu_inst_packet_i_bits_gh_backup; // @[FetchBuffer.scala 85:25]
    end else begin
      fetch_buffer_11_gh_backup <= _GEN_557;
    end
    if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_7 & enq_idxs_7[11]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_11_predict_taken <= io_bpu_inst_packet_i_bits_predict_mask_7; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_6 & enq_idxs_6[11]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_11_predict_taken <= io_bpu_inst_packet_i_bits_predict_mask_6; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_5 & enq_idxs_5[11]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_11_predict_taken <= io_bpu_inst_packet_i_bits_predict_mask_5; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_4 & enq_idxs_4[11]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_11_predict_taken <= io_bpu_inst_packet_i_bits_predict_mask_4; // @[FetchBuffer.scala 85:25]
    end else begin
      fetch_buffer_11_predict_taken <= _GEN_434;
    end
    if (reset) begin // @[FetchBuffer.scala 134:24]
      fetch_buffer_12_inst <= 32'h0; // @[FetchBuffer.scala 17:19]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_7 & enq_idxs_7[12]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_12_inst <= io_bpu_inst_packet_i_bits_data_7; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_6 & enq_idxs_6[12]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_12_inst <= io_bpu_inst_packet_i_bits_data_6; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_5 & enq_idxs_5[12]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_12_inst <= io_bpu_inst_packet_i_bits_data_5; // @[FetchBuffer.scala 85:25]
    end else begin
      fetch_buffer_12_inst <= _GEN_566;
    end
    if (reset) begin // @[FetchBuffer.scala 134:24]
      fetch_buffer_12_inst_addr <= 32'h0; // @[FetchBuffer.scala 18:19]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_7 & enq_idxs_7[12]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_12_inst_addr <= inst_packet_7_inst_addr; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_6 & enq_idxs_6[12]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_12_inst_addr <= inst_packet_6_inst_addr; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_5 & enq_idxs_5[12]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_12_inst_addr <= inst_packet_5_inst_addr; // @[FetchBuffer.scala 85:25]
    end else begin
      fetch_buffer_12_inst_addr <= _GEN_565;
    end
    if (reset) begin // @[FetchBuffer.scala 134:24]
      fetch_buffer_12_gh_backup <= 4'h0; // @[FetchBuffer.scala 19:19]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_7 & enq_idxs_7[12]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_12_gh_backup <= io_bpu_inst_packet_i_bits_gh_backup; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_6 & enq_idxs_6[12]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_12_gh_backup <= io_bpu_inst_packet_i_bits_gh_backup; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_5 & enq_idxs_5[12]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_12_gh_backup <= io_bpu_inst_packet_i_bits_gh_backup; // @[FetchBuffer.scala 85:25]
    end else begin
      fetch_buffer_12_gh_backup <= _GEN_564;
    end
    if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_7 & enq_idxs_7[12]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_12_predict_taken <= io_bpu_inst_packet_i_bits_predict_mask_7; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_6 & enq_idxs_6[12]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_12_predict_taken <= io_bpu_inst_packet_i_bits_predict_mask_6; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_5 & enq_idxs_5[12]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_12_predict_taken <= io_bpu_inst_packet_i_bits_predict_mask_5; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_4 & enq_idxs_4[12]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_12_predict_taken <= io_bpu_inst_packet_i_bits_predict_mask_4; // @[FetchBuffer.scala 85:25]
    end else begin
      fetch_buffer_12_predict_taken <= _GEN_441;
    end
    if (reset) begin // @[FetchBuffer.scala 134:24]
      fetch_buffer_13_inst <= 32'h0; // @[FetchBuffer.scala 17:19]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_7 & enq_idxs_7[13]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_13_inst <= io_bpu_inst_packet_i_bits_data_7; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_6 & enq_idxs_6[13]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_13_inst <= io_bpu_inst_packet_i_bits_data_6; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_5 & enq_idxs_5[13]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_13_inst <= io_bpu_inst_packet_i_bits_data_5; // @[FetchBuffer.scala 85:25]
    end else begin
      fetch_buffer_13_inst <= _GEN_573;
    end
    if (reset) begin // @[FetchBuffer.scala 134:24]
      fetch_buffer_13_inst_addr <= 32'h0; // @[FetchBuffer.scala 18:19]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_7 & enq_idxs_7[13]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_13_inst_addr <= inst_packet_7_inst_addr; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_6 & enq_idxs_6[13]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_13_inst_addr <= inst_packet_6_inst_addr; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_5 & enq_idxs_5[13]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_13_inst_addr <= inst_packet_5_inst_addr; // @[FetchBuffer.scala 85:25]
    end else begin
      fetch_buffer_13_inst_addr <= _GEN_572;
    end
    if (reset) begin // @[FetchBuffer.scala 134:24]
      fetch_buffer_13_gh_backup <= 4'h0; // @[FetchBuffer.scala 19:19]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_7 & enq_idxs_7[13]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_13_gh_backup <= io_bpu_inst_packet_i_bits_gh_backup; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_6 & enq_idxs_6[13]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_13_gh_backup <= io_bpu_inst_packet_i_bits_gh_backup; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_5 & enq_idxs_5[13]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_13_gh_backup <= io_bpu_inst_packet_i_bits_gh_backup; // @[FetchBuffer.scala 85:25]
    end else begin
      fetch_buffer_13_gh_backup <= _GEN_571;
    end
    if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_7 & enq_idxs_7[13]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_13_predict_taken <= io_bpu_inst_packet_i_bits_predict_mask_7; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_6 & enq_idxs_6[13]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_13_predict_taken <= io_bpu_inst_packet_i_bits_predict_mask_6; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_5 & enq_idxs_5[13]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_13_predict_taken <= io_bpu_inst_packet_i_bits_predict_mask_5; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_4 & enq_idxs_4[13]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_13_predict_taken <= io_bpu_inst_packet_i_bits_predict_mask_4; // @[FetchBuffer.scala 85:25]
    end else begin
      fetch_buffer_13_predict_taken <= _GEN_448;
    end
    if (reset) begin // @[FetchBuffer.scala 134:24]
      fetch_buffer_14_inst <= 32'h0; // @[FetchBuffer.scala 17:19]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_7 & enq_idxs_7[14]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_14_inst <= io_bpu_inst_packet_i_bits_data_7; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_6 & enq_idxs_6[14]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_14_inst <= io_bpu_inst_packet_i_bits_data_6; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_5 & enq_idxs_5[14]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_14_inst <= io_bpu_inst_packet_i_bits_data_5; // @[FetchBuffer.scala 85:25]
    end else begin
      fetch_buffer_14_inst <= _GEN_580;
    end
    if (reset) begin // @[FetchBuffer.scala 134:24]
      fetch_buffer_14_inst_addr <= 32'h0; // @[FetchBuffer.scala 18:19]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_7 & enq_idxs_7[14]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_14_inst_addr <= inst_packet_7_inst_addr; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_6 & enq_idxs_6[14]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_14_inst_addr <= inst_packet_6_inst_addr; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_5 & enq_idxs_5[14]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_14_inst_addr <= inst_packet_5_inst_addr; // @[FetchBuffer.scala 85:25]
    end else begin
      fetch_buffer_14_inst_addr <= _GEN_579;
    end
    if (reset) begin // @[FetchBuffer.scala 134:24]
      fetch_buffer_14_gh_backup <= 4'h0; // @[FetchBuffer.scala 19:19]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_7 & enq_idxs_7[14]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_14_gh_backup <= io_bpu_inst_packet_i_bits_gh_backup; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_6 & enq_idxs_6[14]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_14_gh_backup <= io_bpu_inst_packet_i_bits_gh_backup; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_5 & enq_idxs_5[14]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_14_gh_backup <= io_bpu_inst_packet_i_bits_gh_backup; // @[FetchBuffer.scala 85:25]
    end else begin
      fetch_buffer_14_gh_backup <= _GEN_578;
    end
    if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_7 & enq_idxs_7[14]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_14_predict_taken <= io_bpu_inst_packet_i_bits_predict_mask_7; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_6 & enq_idxs_6[14]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_14_predict_taken <= io_bpu_inst_packet_i_bits_predict_mask_6; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_5 & enq_idxs_5[14]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_14_predict_taken <= io_bpu_inst_packet_i_bits_predict_mask_5; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_4 & enq_idxs_4[14]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_14_predict_taken <= io_bpu_inst_packet_i_bits_predict_mask_4; // @[FetchBuffer.scala 85:25]
    end else begin
      fetch_buffer_14_predict_taken <= _GEN_455;
    end
    if (reset) begin // @[FetchBuffer.scala 134:24]
      fetch_buffer_15_inst <= 32'h0; // @[FetchBuffer.scala 17:19]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_7 & enq_idxs_7[15]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_15_inst <= io_bpu_inst_packet_i_bits_data_7; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_6 & enq_idxs_6[15]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_15_inst <= io_bpu_inst_packet_i_bits_data_6; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_5 & enq_idxs_5[15]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_15_inst <= io_bpu_inst_packet_i_bits_data_5; // @[FetchBuffer.scala 85:25]
    end else begin
      fetch_buffer_15_inst <= _GEN_587;
    end
    if (reset) begin // @[FetchBuffer.scala 134:24]
      fetch_buffer_15_inst_addr <= 32'h0; // @[FetchBuffer.scala 18:19]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_7 & enq_idxs_7[15]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_15_inst_addr <= inst_packet_7_inst_addr; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_6 & enq_idxs_6[15]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_15_inst_addr <= inst_packet_6_inst_addr; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_5 & enq_idxs_5[15]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_15_inst_addr <= inst_packet_5_inst_addr; // @[FetchBuffer.scala 85:25]
    end else begin
      fetch_buffer_15_inst_addr <= _GEN_586;
    end
    if (reset) begin // @[FetchBuffer.scala 134:24]
      fetch_buffer_15_gh_backup <= 4'h0; // @[FetchBuffer.scala 19:19]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_7 & enq_idxs_7[15]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_15_gh_backup <= io_bpu_inst_packet_i_bits_gh_backup; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_6 & enq_idxs_6[15]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_15_gh_backup <= io_bpu_inst_packet_i_bits_gh_backup; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_5 & enq_idxs_5[15]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_15_gh_backup <= io_bpu_inst_packet_i_bits_gh_backup; // @[FetchBuffer.scala 85:25]
    end else begin
      fetch_buffer_15_gh_backup <= _GEN_585;
    end
    if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_7 & enq_idxs_7[15]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_15_predict_taken <= io_bpu_inst_packet_i_bits_predict_mask_7; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_6 & enq_idxs_6[15]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_15_predict_taken <= io_bpu_inst_packet_i_bits_predict_mask_6; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_5 & enq_idxs_5[15]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_15_predict_taken <= io_bpu_inst_packet_i_bits_predict_mask_5; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_4 & enq_idxs_4[15]) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_15_predict_taken <= io_bpu_inst_packet_i_bits_predict_mask_4; // @[FetchBuffer.scala 85:25]
    end else begin
      fetch_buffer_15_predict_taken <= _GEN_462;
    end
    if (reset) begin // @[FetchBuffer.scala 134:24]
      fetch_buffer_16_inst <= 32'h0; // @[FetchBuffer.scala 17:19]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_7 & lo_7) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_16_inst <= io_bpu_inst_packet_i_bits_data_7; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_6 & lo_6) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_16_inst <= io_bpu_inst_packet_i_bits_data_6; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_5 & lo_5) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_16_inst <= io_bpu_inst_packet_i_bits_data_5; // @[FetchBuffer.scala 85:25]
    end else begin
      fetch_buffer_16_inst <= _GEN_594;
    end
    if (reset) begin // @[FetchBuffer.scala 134:24]
      fetch_buffer_16_inst_addr <= 32'h0; // @[FetchBuffer.scala 18:19]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_7 & lo_7) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_16_inst_addr <= inst_packet_7_inst_addr; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_6 & lo_6) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_16_inst_addr <= inst_packet_6_inst_addr; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_5 & lo_5) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_16_inst_addr <= inst_packet_5_inst_addr; // @[FetchBuffer.scala 85:25]
    end else begin
      fetch_buffer_16_inst_addr <= _GEN_593;
    end
    if (reset) begin // @[FetchBuffer.scala 134:24]
      fetch_buffer_16_gh_backup <= 4'h0; // @[FetchBuffer.scala 19:19]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_7 & lo_7) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_16_gh_backup <= io_bpu_inst_packet_i_bits_gh_backup; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_6 & lo_6) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_16_gh_backup <= io_bpu_inst_packet_i_bits_gh_backup; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_5 & lo_5) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_16_gh_backup <= io_bpu_inst_packet_i_bits_gh_backup; // @[FetchBuffer.scala 85:25]
    end else begin
      fetch_buffer_16_gh_backup <= _GEN_592;
    end
    if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_7 & lo_7) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_16_predict_taken <= io_bpu_inst_packet_i_bits_predict_mask_7; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_6 & lo_6) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_16_predict_taken <= io_bpu_inst_packet_i_bits_predict_mask_6; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_5 & lo_5) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_16_predict_taken <= io_bpu_inst_packet_i_bits_predict_mask_5; // @[FetchBuffer.scala 85:25]
    end else if (do_enq & io_bpu_inst_packet_i_bits_valid_mask_4 & lo_4) begin // @[FetchBuffer.scala 84:65]
      fetch_buffer_16_predict_taken <= io_bpu_inst_packet_i_bits_predict_mask_4; // @[FetchBuffer.scala 85:25]
    end else begin
      fetch_buffer_16_predict_taken <= _GEN_469;
    end
    if (reset) begin // @[FetchBuffer.scala 51:29]
      deq_idxs_0 <= 17'h1; // @[FetchBuffer.scala 51:29]
    end else if (io_clear_i) begin // @[FetchBuffer.scala 125:20]
      deq_idxs_0 <= 17'h1; // @[FetchBuffer.scala 127:10]
    end else if (io_fb_resp_deq_valid_1) begin // @[FetchBuffer.scala 111:20]
      deq_idxs_0 <= _T_459;
    end else if (io_fb_resp_deq_valid_0) begin // @[FetchBuffer.scala 111:20]
      deq_idxs_0 <= deq_idxs_1;
    end
    if (reset) begin // @[FetchBuffer.scala 52:29]
      tail <= 17'h1; // @[FetchBuffer.scala 52:29]
    end else if (io_clear_i) begin // @[FetchBuffer.scala 125:20]
      tail <= 17'h1; // @[FetchBuffer.scala 126:10]
    end else if (do_enq) begin // @[FetchBuffer.scala 89:16]
      if (io_bpu_inst_packet_i_bits_valid_mask_7) begin // @[FetchBuffer.scala 68:18]
        tail <= _T_14;
      end else begin
        tail <= enq_idxs_7;
      end
    end
    if (reset) begin // @[FetchBuffer.scala 53:29]
      maybe_full <= 1'h0; // @[FetchBuffer.scala 53:29]
    end else if (io_clear_i) begin // @[FetchBuffer.scala 125:20]
      maybe_full <= 1'h0; // @[FetchBuffer.scala 128:16]
    end else begin
      maybe_full <= _GEN_1193;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  fetch_buffer_0_inst = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  fetch_buffer_0_inst_addr = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  fetch_buffer_0_gh_backup = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  fetch_buffer_0_predict_taken = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  fetch_buffer_1_inst = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  fetch_buffer_1_inst_addr = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  fetch_buffer_1_gh_backup = _RAND_6[3:0];
  _RAND_7 = {1{`RANDOM}};
  fetch_buffer_1_predict_taken = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  fetch_buffer_2_inst = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  fetch_buffer_2_inst_addr = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  fetch_buffer_2_gh_backup = _RAND_10[3:0];
  _RAND_11 = {1{`RANDOM}};
  fetch_buffer_2_predict_taken = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  fetch_buffer_3_inst = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  fetch_buffer_3_inst_addr = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  fetch_buffer_3_gh_backup = _RAND_14[3:0];
  _RAND_15 = {1{`RANDOM}};
  fetch_buffer_3_predict_taken = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  fetch_buffer_4_inst = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  fetch_buffer_4_inst_addr = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  fetch_buffer_4_gh_backup = _RAND_18[3:0];
  _RAND_19 = {1{`RANDOM}};
  fetch_buffer_4_predict_taken = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  fetch_buffer_5_inst = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  fetch_buffer_5_inst_addr = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  fetch_buffer_5_gh_backup = _RAND_22[3:0];
  _RAND_23 = {1{`RANDOM}};
  fetch_buffer_5_predict_taken = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  fetch_buffer_6_inst = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  fetch_buffer_6_inst_addr = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  fetch_buffer_6_gh_backup = _RAND_26[3:0];
  _RAND_27 = {1{`RANDOM}};
  fetch_buffer_6_predict_taken = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  fetch_buffer_7_inst = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  fetch_buffer_7_inst_addr = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  fetch_buffer_7_gh_backup = _RAND_30[3:0];
  _RAND_31 = {1{`RANDOM}};
  fetch_buffer_7_predict_taken = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  fetch_buffer_8_inst = _RAND_32[31:0];
  _RAND_33 = {1{`RANDOM}};
  fetch_buffer_8_inst_addr = _RAND_33[31:0];
  _RAND_34 = {1{`RANDOM}};
  fetch_buffer_8_gh_backup = _RAND_34[3:0];
  _RAND_35 = {1{`RANDOM}};
  fetch_buffer_8_predict_taken = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  fetch_buffer_9_inst = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  fetch_buffer_9_inst_addr = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  fetch_buffer_9_gh_backup = _RAND_38[3:0];
  _RAND_39 = {1{`RANDOM}};
  fetch_buffer_9_predict_taken = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  fetch_buffer_10_inst = _RAND_40[31:0];
  _RAND_41 = {1{`RANDOM}};
  fetch_buffer_10_inst_addr = _RAND_41[31:0];
  _RAND_42 = {1{`RANDOM}};
  fetch_buffer_10_gh_backup = _RAND_42[3:0];
  _RAND_43 = {1{`RANDOM}};
  fetch_buffer_10_predict_taken = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  fetch_buffer_11_inst = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  fetch_buffer_11_inst_addr = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  fetch_buffer_11_gh_backup = _RAND_46[3:0];
  _RAND_47 = {1{`RANDOM}};
  fetch_buffer_11_predict_taken = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  fetch_buffer_12_inst = _RAND_48[31:0];
  _RAND_49 = {1{`RANDOM}};
  fetch_buffer_12_inst_addr = _RAND_49[31:0];
  _RAND_50 = {1{`RANDOM}};
  fetch_buffer_12_gh_backup = _RAND_50[3:0];
  _RAND_51 = {1{`RANDOM}};
  fetch_buffer_12_predict_taken = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  fetch_buffer_13_inst = _RAND_52[31:0];
  _RAND_53 = {1{`RANDOM}};
  fetch_buffer_13_inst_addr = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  fetch_buffer_13_gh_backup = _RAND_54[3:0];
  _RAND_55 = {1{`RANDOM}};
  fetch_buffer_13_predict_taken = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  fetch_buffer_14_inst = _RAND_56[31:0];
  _RAND_57 = {1{`RANDOM}};
  fetch_buffer_14_inst_addr = _RAND_57[31:0];
  _RAND_58 = {1{`RANDOM}};
  fetch_buffer_14_gh_backup = _RAND_58[3:0];
  _RAND_59 = {1{`RANDOM}};
  fetch_buffer_14_predict_taken = _RAND_59[0:0];
  _RAND_60 = {1{`RANDOM}};
  fetch_buffer_15_inst = _RAND_60[31:0];
  _RAND_61 = {1{`RANDOM}};
  fetch_buffer_15_inst_addr = _RAND_61[31:0];
  _RAND_62 = {1{`RANDOM}};
  fetch_buffer_15_gh_backup = _RAND_62[3:0];
  _RAND_63 = {1{`RANDOM}};
  fetch_buffer_15_predict_taken = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  fetch_buffer_16_inst = _RAND_64[31:0];
  _RAND_65 = {1{`RANDOM}};
  fetch_buffer_16_inst_addr = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  fetch_buffer_16_gh_backup = _RAND_66[3:0];
  _RAND_67 = {1{`RANDOM}};
  fetch_buffer_16_predict_taken = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  deq_idxs_0 = _RAND_68[16:0];
  _RAND_69 = {1{`RANDOM}};
  tail = _RAND_69[16:0];
  _RAND_70 = {1{`RANDOM}};
  maybe_full = _RAND_70[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Ifu(
  input          clock,
  input          reset,
  input          io_ex_branch_info_i_valid,
  input  [31:0]  io_ex_branch_info_i_bits_target_addr,
  input  [31:0]  io_ex_branch_info_i_bits_inst_addr,
  input  [3:0]   io_ex_branch_info_i_bits_gh_update,
  input          io_ex_branch_info_i_bits_is_branch,
  input          io_ex_branch_info_i_bits_is_taken,
  input          io_ex_branch_info_i_bits_predict_miss,
  output         io_fb_inst_bank_o_valid,
  output [31:0]  io_fb_inst_bank_o_bits_data_0_inst,
  output [31:0]  io_fb_inst_bank_o_bits_data_0_inst_addr,
  output [3:0]   io_fb_inst_bank_o_bits_data_0_gh_backup,
  output         io_fb_inst_bank_o_bits_data_0_is_valid,
  output         io_fb_inst_bank_o_bits_data_0_predict_taken,
  output [31:0]  io_fb_inst_bank_o_bits_data_1_inst,
  output [31:0]  io_fb_inst_bank_o_bits_data_1_inst_addr,
  output [3:0]   io_fb_inst_bank_o_bits_data_1_gh_backup,
  output         io_fb_inst_bank_o_bits_data_1_is_valid,
  output         io_fb_inst_bank_o_bits_data_1_predict_taken,
  input          io_fb_resp_deq_valid_0,
  input          io_fb_resp_deq_valid_1,
  input          io_icache_io_read_req_ready,
  output         io_icache_io_read_req_valid,
  output [31:0]  io_icache_io_read_req_bits_addr,
  input  [255:0] io_icache_io_read_resp_bits_data,
  output         io_icache_debug_state,
  output         io_icache_debug_hit_cache,
  output         io_icache_debug_cache_we,
  output [19:0]  io_icache_debug_cache_read_tag,
  output         io_icache_debug_icache_req_valid,
  output [31:0]  io_icache_debug_icache_req_bits_addr,
  output [7:0]   io_bpu_debug_branch_mask,
  output [7:0]   io_bpu_debug_fetched_mask,
  output [7:0]   io_bpu_debug_predict_branch,
  output [31:0]  io_bpu_debug_predict_addr,
  output         io_bpu_debug_is_taken,
  output         io_bpu_debug_take_delay,
  output [31:0]  io_bpu_debug_inst_packet_0,
  output [31:0]  io_bpu_debug_inst_packet_1,
  output [31:0]  io_bpu_debug_inst_packet_2,
  output [31:0]  io_bpu_debug_inst_packet_3,
  output [31:0]  io_bpu_debug_inst_packet_4,
  output [31:0]  io_bpu_debug_inst_packet_5,
  output [31:0]  io_bpu_debug_inst_packet_6,
  output [31:0]  io_bpu_debug_inst_packet_7
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  bpu_clock; // @[Ifu.scala 19:28]
  wire  bpu_reset; // @[Ifu.scala 19:28]
  wire  bpu_io_inst_packet_i_valid; // @[Ifu.scala 19:28]
  wire [31:0] bpu_io_inst_packet_i_bits_data_0; // @[Ifu.scala 19:28]
  wire [31:0] bpu_io_inst_packet_i_bits_data_1; // @[Ifu.scala 19:28]
  wire [31:0] bpu_io_inst_packet_i_bits_data_2; // @[Ifu.scala 19:28]
  wire [31:0] bpu_io_inst_packet_i_bits_data_3; // @[Ifu.scala 19:28]
  wire [31:0] bpu_io_inst_packet_i_bits_data_4; // @[Ifu.scala 19:28]
  wire [31:0] bpu_io_inst_packet_i_bits_data_5; // @[Ifu.scala 19:28]
  wire [31:0] bpu_io_inst_packet_i_bits_data_6; // @[Ifu.scala 19:28]
  wire [31:0] bpu_io_inst_packet_i_bits_data_7; // @[Ifu.scala 19:28]
  wire [31:0] bpu_io_inst_packet_i_bits_addr; // @[Ifu.scala 19:28]
  wire  bpu_io_resp_o_valid; // @[Ifu.scala 19:28]
  wire [31:0] bpu_io_resp_o_bits_predict_addr; // @[Ifu.scala 19:28]
  wire  bpu_io_resp_o_bits_is_taken; // @[Ifu.scala 19:28]
  wire  bpu_io_resp_o_bits_take_delay; // @[Ifu.scala 19:28]
  wire  bpu_io_bpu_inst_packet_o_ready; // @[Ifu.scala 19:28]
  wire  bpu_io_bpu_inst_packet_o_valid; // @[Ifu.scala 19:28]
  wire [31:0] bpu_io_bpu_inst_packet_o_bits_data_0; // @[Ifu.scala 19:28]
  wire [31:0] bpu_io_bpu_inst_packet_o_bits_data_1; // @[Ifu.scala 19:28]
  wire [31:0] bpu_io_bpu_inst_packet_o_bits_data_2; // @[Ifu.scala 19:28]
  wire [31:0] bpu_io_bpu_inst_packet_o_bits_data_3; // @[Ifu.scala 19:28]
  wire [31:0] bpu_io_bpu_inst_packet_o_bits_data_4; // @[Ifu.scala 19:28]
  wire [31:0] bpu_io_bpu_inst_packet_o_bits_data_5; // @[Ifu.scala 19:28]
  wire [31:0] bpu_io_bpu_inst_packet_o_bits_data_6; // @[Ifu.scala 19:28]
  wire [31:0] bpu_io_bpu_inst_packet_o_bits_data_7; // @[Ifu.scala 19:28]
  wire [31:0] bpu_io_bpu_inst_packet_o_bits_addr; // @[Ifu.scala 19:28]
  wire [3:0] bpu_io_bpu_inst_packet_o_bits_gh_backup; // @[Ifu.scala 19:28]
  wire  bpu_io_bpu_inst_packet_o_bits_valid_mask_0; // @[Ifu.scala 19:28]
  wire  bpu_io_bpu_inst_packet_o_bits_valid_mask_1; // @[Ifu.scala 19:28]
  wire  bpu_io_bpu_inst_packet_o_bits_valid_mask_2; // @[Ifu.scala 19:28]
  wire  bpu_io_bpu_inst_packet_o_bits_valid_mask_3; // @[Ifu.scala 19:28]
  wire  bpu_io_bpu_inst_packet_o_bits_valid_mask_4; // @[Ifu.scala 19:28]
  wire  bpu_io_bpu_inst_packet_o_bits_valid_mask_5; // @[Ifu.scala 19:28]
  wire  bpu_io_bpu_inst_packet_o_bits_valid_mask_6; // @[Ifu.scala 19:28]
  wire  bpu_io_bpu_inst_packet_o_bits_valid_mask_7; // @[Ifu.scala 19:28]
  wire  bpu_io_bpu_inst_packet_o_bits_predict_mask_0; // @[Ifu.scala 19:28]
  wire  bpu_io_bpu_inst_packet_o_bits_predict_mask_1; // @[Ifu.scala 19:28]
  wire  bpu_io_bpu_inst_packet_o_bits_predict_mask_2; // @[Ifu.scala 19:28]
  wire  bpu_io_bpu_inst_packet_o_bits_predict_mask_3; // @[Ifu.scala 19:28]
  wire  bpu_io_bpu_inst_packet_o_bits_predict_mask_4; // @[Ifu.scala 19:28]
  wire  bpu_io_bpu_inst_packet_o_bits_predict_mask_5; // @[Ifu.scala 19:28]
  wire  bpu_io_bpu_inst_packet_o_bits_predict_mask_6; // @[Ifu.scala 19:28]
  wire  bpu_io_bpu_inst_packet_o_bits_predict_mask_7; // @[Ifu.scala 19:28]
  wire  bpu_io_branch_info_i_valid; // @[Ifu.scala 19:28]
  wire [31:0] bpu_io_branch_info_i_bits_inst_addr; // @[Ifu.scala 19:28]
  wire [3:0] bpu_io_branch_info_i_bits_gh_update; // @[Ifu.scala 19:28]
  wire  bpu_io_branch_info_i_bits_is_branch; // @[Ifu.scala 19:28]
  wire  bpu_io_branch_info_i_bits_is_taken; // @[Ifu.scala 19:28]
  wire  bpu_io_branch_info_i_bits_predict_miss; // @[Ifu.scala 19:28]
  wire  bpu_io_is_delay; // @[Ifu.scala 19:28]
  wire  bpu_io_need_flush; // @[Ifu.scala 19:28]
  wire [7:0] bpu_io_bpu_debug_branch_mask; // @[Ifu.scala 19:28]
  wire [7:0] bpu_io_bpu_debug_fetched_mask; // @[Ifu.scala 19:28]
  wire [7:0] bpu_io_bpu_debug_predict_branch; // @[Ifu.scala 19:28]
  wire [31:0] bpu_io_bpu_debug_predict_addr; // @[Ifu.scala 19:28]
  wire  bpu_io_bpu_debug_is_taken; // @[Ifu.scala 19:28]
  wire  bpu_io_bpu_debug_take_delay; // @[Ifu.scala 19:28]
  wire [31:0] bpu_io_bpu_debug_inst_packet_0; // @[Ifu.scala 19:28]
  wire [31:0] bpu_io_bpu_debug_inst_packet_1; // @[Ifu.scala 19:28]
  wire [31:0] bpu_io_bpu_debug_inst_packet_2; // @[Ifu.scala 19:28]
  wire [31:0] bpu_io_bpu_debug_inst_packet_3; // @[Ifu.scala 19:28]
  wire [31:0] bpu_io_bpu_debug_inst_packet_4; // @[Ifu.scala 19:28]
  wire [31:0] bpu_io_bpu_debug_inst_packet_5; // @[Ifu.scala 19:28]
  wire [31:0] bpu_io_bpu_debug_inst_packet_6; // @[Ifu.scala 19:28]
  wire [31:0] bpu_io_bpu_debug_inst_packet_7; // @[Ifu.scala 19:28]
  wire  icache_clock; // @[Ifu.scala 20:28]
  wire  icache_reset; // @[Ifu.scala 20:28]
  wire  icache_io_icache_req_ready; // @[Ifu.scala 20:28]
  wire  icache_io_icache_req_valid; // @[Ifu.scala 20:28]
  wire [31:0] icache_io_icache_req_bits_addr; // @[Ifu.scala 20:28]
  wire  icache_io_icache_resp_valid; // @[Ifu.scala 20:28]
  wire [31:0] icache_io_icache_resp_bits_data_0; // @[Ifu.scala 20:28]
  wire [31:0] icache_io_icache_resp_bits_data_1; // @[Ifu.scala 20:28]
  wire [31:0] icache_io_icache_resp_bits_data_2; // @[Ifu.scala 20:28]
  wire [31:0] icache_io_icache_resp_bits_data_3; // @[Ifu.scala 20:28]
  wire [31:0] icache_io_icache_resp_bits_data_4; // @[Ifu.scala 20:28]
  wire [31:0] icache_io_icache_resp_bits_data_5; // @[Ifu.scala 20:28]
  wire [31:0] icache_io_icache_resp_bits_data_6; // @[Ifu.scala 20:28]
  wire [31:0] icache_io_icache_resp_bits_data_7; // @[Ifu.scala 20:28]
  wire [31:0] icache_io_icache_resp_bits_addr; // @[Ifu.scala 20:28]
  wire  icache_io_io_read_req_ready; // @[Ifu.scala 20:28]
  wire  icache_io_io_read_req_valid; // @[Ifu.scala 20:28]
  wire [31:0] icache_io_io_read_req_bits_addr; // @[Ifu.scala 20:28]
  wire [255:0] icache_io_io_read_resp_bits_data; // @[Ifu.scala 20:28]
  wire  icache_io_icache_debug_state; // @[Ifu.scala 20:28]
  wire  icache_io_icache_debug_hit_cache; // @[Ifu.scala 20:28]
  wire  icache_io_icache_debug_cache_we; // @[Ifu.scala 20:28]
  wire [19:0] icache_io_icache_debug_cache_read_tag; // @[Ifu.scala 20:28]
  wire  icache_io_icache_debug_icache_req_valid; // @[Ifu.scala 20:28]
  wire [31:0] icache_io_icache_debug_icache_req_bits_addr; // @[Ifu.scala 20:28]
  wire  fetch_buffer_clock; // @[Ifu.scala 21:28]
  wire  fetch_buffer_reset; // @[Ifu.scala 21:28]
  wire  fetch_buffer_io_bpu_inst_packet_i_ready; // @[Ifu.scala 21:28]
  wire  fetch_buffer_io_bpu_inst_packet_i_valid; // @[Ifu.scala 21:28]
  wire [31:0] fetch_buffer_io_bpu_inst_packet_i_bits_data_0; // @[Ifu.scala 21:28]
  wire [31:0] fetch_buffer_io_bpu_inst_packet_i_bits_data_1; // @[Ifu.scala 21:28]
  wire [31:0] fetch_buffer_io_bpu_inst_packet_i_bits_data_2; // @[Ifu.scala 21:28]
  wire [31:0] fetch_buffer_io_bpu_inst_packet_i_bits_data_3; // @[Ifu.scala 21:28]
  wire [31:0] fetch_buffer_io_bpu_inst_packet_i_bits_data_4; // @[Ifu.scala 21:28]
  wire [31:0] fetch_buffer_io_bpu_inst_packet_i_bits_data_5; // @[Ifu.scala 21:28]
  wire [31:0] fetch_buffer_io_bpu_inst_packet_i_bits_data_6; // @[Ifu.scala 21:28]
  wire [31:0] fetch_buffer_io_bpu_inst_packet_i_bits_data_7; // @[Ifu.scala 21:28]
  wire [31:0] fetch_buffer_io_bpu_inst_packet_i_bits_addr; // @[Ifu.scala 21:28]
  wire [3:0] fetch_buffer_io_bpu_inst_packet_i_bits_gh_backup; // @[Ifu.scala 21:28]
  wire  fetch_buffer_io_bpu_inst_packet_i_bits_valid_mask_0; // @[Ifu.scala 21:28]
  wire  fetch_buffer_io_bpu_inst_packet_i_bits_valid_mask_1; // @[Ifu.scala 21:28]
  wire  fetch_buffer_io_bpu_inst_packet_i_bits_valid_mask_2; // @[Ifu.scala 21:28]
  wire  fetch_buffer_io_bpu_inst_packet_i_bits_valid_mask_3; // @[Ifu.scala 21:28]
  wire  fetch_buffer_io_bpu_inst_packet_i_bits_valid_mask_4; // @[Ifu.scala 21:28]
  wire  fetch_buffer_io_bpu_inst_packet_i_bits_valid_mask_5; // @[Ifu.scala 21:28]
  wire  fetch_buffer_io_bpu_inst_packet_i_bits_valid_mask_6; // @[Ifu.scala 21:28]
  wire  fetch_buffer_io_bpu_inst_packet_i_bits_valid_mask_7; // @[Ifu.scala 21:28]
  wire  fetch_buffer_io_bpu_inst_packet_i_bits_predict_mask_0; // @[Ifu.scala 21:28]
  wire  fetch_buffer_io_bpu_inst_packet_i_bits_predict_mask_1; // @[Ifu.scala 21:28]
  wire  fetch_buffer_io_bpu_inst_packet_i_bits_predict_mask_2; // @[Ifu.scala 21:28]
  wire  fetch_buffer_io_bpu_inst_packet_i_bits_predict_mask_3; // @[Ifu.scala 21:28]
  wire  fetch_buffer_io_bpu_inst_packet_i_bits_predict_mask_4; // @[Ifu.scala 21:28]
  wire  fetch_buffer_io_bpu_inst_packet_i_bits_predict_mask_5; // @[Ifu.scala 21:28]
  wire  fetch_buffer_io_bpu_inst_packet_i_bits_predict_mask_6; // @[Ifu.scala 21:28]
  wire  fetch_buffer_io_bpu_inst_packet_i_bits_predict_mask_7; // @[Ifu.scala 21:28]
  wire  fetch_buffer_io_inst_bank_valid; // @[Ifu.scala 21:28]
  wire [31:0] fetch_buffer_io_inst_bank_bits_data_0_inst; // @[Ifu.scala 21:28]
  wire [31:0] fetch_buffer_io_inst_bank_bits_data_0_inst_addr; // @[Ifu.scala 21:28]
  wire [3:0] fetch_buffer_io_inst_bank_bits_data_0_gh_backup; // @[Ifu.scala 21:28]
  wire  fetch_buffer_io_inst_bank_bits_data_0_is_valid; // @[Ifu.scala 21:28]
  wire  fetch_buffer_io_inst_bank_bits_data_0_predict_taken; // @[Ifu.scala 21:28]
  wire [31:0] fetch_buffer_io_inst_bank_bits_data_1_inst; // @[Ifu.scala 21:28]
  wire [31:0] fetch_buffer_io_inst_bank_bits_data_1_inst_addr; // @[Ifu.scala 21:28]
  wire [3:0] fetch_buffer_io_inst_bank_bits_data_1_gh_backup; // @[Ifu.scala 21:28]
  wire  fetch_buffer_io_inst_bank_bits_data_1_is_valid; // @[Ifu.scala 21:28]
  wire  fetch_buffer_io_inst_bank_bits_data_1_predict_taken; // @[Ifu.scala 21:28]
  wire  fetch_buffer_io_fb_resp_deq_valid_0; // @[Ifu.scala 21:28]
  wire  fetch_buffer_io_fb_resp_deq_valid_1; // @[Ifu.scala 21:28]
  wire  fetch_buffer_io_clear_i; // @[Ifu.scala 21:28]
  reg [31:0] pc; // @[Ifu.scala 23:30]
  wire [26:0] no_taken_addr_hi = pc[31:5] + 27'h1; // @[Ifu.scala 24:56]
  wire [31:0] no_taken_addr = {no_taken_addr_hi,5'h0}; // @[Cat.scala 30:58]
  wire  stop_fetch = ~fetch_buffer_io_bpu_inst_packet_i_ready | ~icache_io_icache_req_ready | ~bpu_io_resp_o_valid; // @[Ifu.scala 25:92]
  wire  redirect = io_ex_branch_info_i_valid & io_ex_branch_info_i_bits_predict_miss; // @[Ifu.scala 26:44]
  reg  taking_delay; // @[Ifu.scala 28:34]
  reg [31:0] delay_target_addr; // @[Ifu.scala 29:34]
  wire [31:0] _GEN_0 = bpu_io_resp_o_bits_is_taken ? bpu_io_resp_o_bits_predict_addr : no_taken_addr; // @[Ifu.scala 43:43 Ifu.scala 44:8 Ifu.scala 46:8]
  wire [31:0] _GEN_1 = bpu_io_resp_o_bits_take_delay ? no_taken_addr : _GEN_0; // @[Ifu.scala 39:45 Ifu.scala 40:8]
  wire  _GEN_2 = bpu_io_resp_o_bits_take_delay | taking_delay; // @[Ifu.scala 39:45 Ifu.scala 41:18 Ifu.scala 28:34]
  wire [31:0] _GEN_3 = bpu_io_resp_o_bits_take_delay ? bpu_io_resp_o_bits_predict_addr : delay_target_addr; // @[Ifu.scala 39:45 Ifu.scala 42:23 Ifu.scala 29:34]
  BPU bpu ( // @[Ifu.scala 19:28]
    .clock(bpu_clock),
    .reset(bpu_reset),
    .io_inst_packet_i_valid(bpu_io_inst_packet_i_valid),
    .io_inst_packet_i_bits_data_0(bpu_io_inst_packet_i_bits_data_0),
    .io_inst_packet_i_bits_data_1(bpu_io_inst_packet_i_bits_data_1),
    .io_inst_packet_i_bits_data_2(bpu_io_inst_packet_i_bits_data_2),
    .io_inst_packet_i_bits_data_3(bpu_io_inst_packet_i_bits_data_3),
    .io_inst_packet_i_bits_data_4(bpu_io_inst_packet_i_bits_data_4),
    .io_inst_packet_i_bits_data_5(bpu_io_inst_packet_i_bits_data_5),
    .io_inst_packet_i_bits_data_6(bpu_io_inst_packet_i_bits_data_6),
    .io_inst_packet_i_bits_data_7(bpu_io_inst_packet_i_bits_data_7),
    .io_inst_packet_i_bits_addr(bpu_io_inst_packet_i_bits_addr),
    .io_resp_o_valid(bpu_io_resp_o_valid),
    .io_resp_o_bits_predict_addr(bpu_io_resp_o_bits_predict_addr),
    .io_resp_o_bits_is_taken(bpu_io_resp_o_bits_is_taken),
    .io_resp_o_bits_take_delay(bpu_io_resp_o_bits_take_delay),
    .io_bpu_inst_packet_o_ready(bpu_io_bpu_inst_packet_o_ready),
    .io_bpu_inst_packet_o_valid(bpu_io_bpu_inst_packet_o_valid),
    .io_bpu_inst_packet_o_bits_data_0(bpu_io_bpu_inst_packet_o_bits_data_0),
    .io_bpu_inst_packet_o_bits_data_1(bpu_io_bpu_inst_packet_o_bits_data_1),
    .io_bpu_inst_packet_o_bits_data_2(bpu_io_bpu_inst_packet_o_bits_data_2),
    .io_bpu_inst_packet_o_bits_data_3(bpu_io_bpu_inst_packet_o_bits_data_3),
    .io_bpu_inst_packet_o_bits_data_4(bpu_io_bpu_inst_packet_o_bits_data_4),
    .io_bpu_inst_packet_o_bits_data_5(bpu_io_bpu_inst_packet_o_bits_data_5),
    .io_bpu_inst_packet_o_bits_data_6(bpu_io_bpu_inst_packet_o_bits_data_6),
    .io_bpu_inst_packet_o_bits_data_7(bpu_io_bpu_inst_packet_o_bits_data_7),
    .io_bpu_inst_packet_o_bits_addr(bpu_io_bpu_inst_packet_o_bits_addr),
    .io_bpu_inst_packet_o_bits_gh_backup(bpu_io_bpu_inst_packet_o_bits_gh_backup),
    .io_bpu_inst_packet_o_bits_valid_mask_0(bpu_io_bpu_inst_packet_o_bits_valid_mask_0),
    .io_bpu_inst_packet_o_bits_valid_mask_1(bpu_io_bpu_inst_packet_o_bits_valid_mask_1),
    .io_bpu_inst_packet_o_bits_valid_mask_2(bpu_io_bpu_inst_packet_o_bits_valid_mask_2),
    .io_bpu_inst_packet_o_bits_valid_mask_3(bpu_io_bpu_inst_packet_o_bits_valid_mask_3),
    .io_bpu_inst_packet_o_bits_valid_mask_4(bpu_io_bpu_inst_packet_o_bits_valid_mask_4),
    .io_bpu_inst_packet_o_bits_valid_mask_5(bpu_io_bpu_inst_packet_o_bits_valid_mask_5),
    .io_bpu_inst_packet_o_bits_valid_mask_6(bpu_io_bpu_inst_packet_o_bits_valid_mask_6),
    .io_bpu_inst_packet_o_bits_valid_mask_7(bpu_io_bpu_inst_packet_o_bits_valid_mask_7),
    .io_bpu_inst_packet_o_bits_predict_mask_0(bpu_io_bpu_inst_packet_o_bits_predict_mask_0),
    .io_bpu_inst_packet_o_bits_predict_mask_1(bpu_io_bpu_inst_packet_o_bits_predict_mask_1),
    .io_bpu_inst_packet_o_bits_predict_mask_2(bpu_io_bpu_inst_packet_o_bits_predict_mask_2),
    .io_bpu_inst_packet_o_bits_predict_mask_3(bpu_io_bpu_inst_packet_o_bits_predict_mask_3),
    .io_bpu_inst_packet_o_bits_predict_mask_4(bpu_io_bpu_inst_packet_o_bits_predict_mask_4),
    .io_bpu_inst_packet_o_bits_predict_mask_5(bpu_io_bpu_inst_packet_o_bits_predict_mask_5),
    .io_bpu_inst_packet_o_bits_predict_mask_6(bpu_io_bpu_inst_packet_o_bits_predict_mask_6),
    .io_bpu_inst_packet_o_bits_predict_mask_7(bpu_io_bpu_inst_packet_o_bits_predict_mask_7),
    .io_branch_info_i_valid(bpu_io_branch_info_i_valid),
    .io_branch_info_i_bits_inst_addr(bpu_io_branch_info_i_bits_inst_addr),
    .io_branch_info_i_bits_gh_update(bpu_io_branch_info_i_bits_gh_update),
    .io_branch_info_i_bits_is_branch(bpu_io_branch_info_i_bits_is_branch),
    .io_branch_info_i_bits_is_taken(bpu_io_branch_info_i_bits_is_taken),
    .io_branch_info_i_bits_predict_miss(bpu_io_branch_info_i_bits_predict_miss),
    .io_is_delay(bpu_io_is_delay),
    .io_need_flush(bpu_io_need_flush),
    .io_bpu_debug_branch_mask(bpu_io_bpu_debug_branch_mask),
    .io_bpu_debug_fetched_mask(bpu_io_bpu_debug_fetched_mask),
    .io_bpu_debug_predict_branch(bpu_io_bpu_debug_predict_branch),
    .io_bpu_debug_predict_addr(bpu_io_bpu_debug_predict_addr),
    .io_bpu_debug_is_taken(bpu_io_bpu_debug_is_taken),
    .io_bpu_debug_take_delay(bpu_io_bpu_debug_take_delay),
    .io_bpu_debug_inst_packet_0(bpu_io_bpu_debug_inst_packet_0),
    .io_bpu_debug_inst_packet_1(bpu_io_bpu_debug_inst_packet_1),
    .io_bpu_debug_inst_packet_2(bpu_io_bpu_debug_inst_packet_2),
    .io_bpu_debug_inst_packet_3(bpu_io_bpu_debug_inst_packet_3),
    .io_bpu_debug_inst_packet_4(bpu_io_bpu_debug_inst_packet_4),
    .io_bpu_debug_inst_packet_5(bpu_io_bpu_debug_inst_packet_5),
    .io_bpu_debug_inst_packet_6(bpu_io_bpu_debug_inst_packet_6),
    .io_bpu_debug_inst_packet_7(bpu_io_bpu_debug_inst_packet_7)
  );
  ICache icache ( // @[Ifu.scala 20:28]
    .clock(icache_clock),
    .reset(icache_reset),
    .io_icache_req_ready(icache_io_icache_req_ready),
    .io_icache_req_valid(icache_io_icache_req_valid),
    .io_icache_req_bits_addr(icache_io_icache_req_bits_addr),
    .io_icache_resp_valid(icache_io_icache_resp_valid),
    .io_icache_resp_bits_data_0(icache_io_icache_resp_bits_data_0),
    .io_icache_resp_bits_data_1(icache_io_icache_resp_bits_data_1),
    .io_icache_resp_bits_data_2(icache_io_icache_resp_bits_data_2),
    .io_icache_resp_bits_data_3(icache_io_icache_resp_bits_data_3),
    .io_icache_resp_bits_data_4(icache_io_icache_resp_bits_data_4),
    .io_icache_resp_bits_data_5(icache_io_icache_resp_bits_data_5),
    .io_icache_resp_bits_data_6(icache_io_icache_resp_bits_data_6),
    .io_icache_resp_bits_data_7(icache_io_icache_resp_bits_data_7),
    .io_icache_resp_bits_addr(icache_io_icache_resp_bits_addr),
    .io_io_read_req_ready(icache_io_io_read_req_ready),
    .io_io_read_req_valid(icache_io_io_read_req_valid),
    .io_io_read_req_bits_addr(icache_io_io_read_req_bits_addr),
    .io_io_read_resp_bits_data(icache_io_io_read_resp_bits_data),
    .io_icache_debug_state(icache_io_icache_debug_state),
    .io_icache_debug_hit_cache(icache_io_icache_debug_hit_cache),
    .io_icache_debug_cache_we(icache_io_icache_debug_cache_we),
    .io_icache_debug_cache_read_tag(icache_io_icache_debug_cache_read_tag),
    .io_icache_debug_icache_req_valid(icache_io_icache_debug_icache_req_valid),
    .io_icache_debug_icache_req_bits_addr(icache_io_icache_debug_icache_req_bits_addr)
  );
  FetchBuffer fetch_buffer ( // @[Ifu.scala 21:28]
    .clock(fetch_buffer_clock),
    .reset(fetch_buffer_reset),
    .io_bpu_inst_packet_i_ready(fetch_buffer_io_bpu_inst_packet_i_ready),
    .io_bpu_inst_packet_i_valid(fetch_buffer_io_bpu_inst_packet_i_valid),
    .io_bpu_inst_packet_i_bits_data_0(fetch_buffer_io_bpu_inst_packet_i_bits_data_0),
    .io_bpu_inst_packet_i_bits_data_1(fetch_buffer_io_bpu_inst_packet_i_bits_data_1),
    .io_bpu_inst_packet_i_bits_data_2(fetch_buffer_io_bpu_inst_packet_i_bits_data_2),
    .io_bpu_inst_packet_i_bits_data_3(fetch_buffer_io_bpu_inst_packet_i_bits_data_3),
    .io_bpu_inst_packet_i_bits_data_4(fetch_buffer_io_bpu_inst_packet_i_bits_data_4),
    .io_bpu_inst_packet_i_bits_data_5(fetch_buffer_io_bpu_inst_packet_i_bits_data_5),
    .io_bpu_inst_packet_i_bits_data_6(fetch_buffer_io_bpu_inst_packet_i_bits_data_6),
    .io_bpu_inst_packet_i_bits_data_7(fetch_buffer_io_bpu_inst_packet_i_bits_data_7),
    .io_bpu_inst_packet_i_bits_addr(fetch_buffer_io_bpu_inst_packet_i_bits_addr),
    .io_bpu_inst_packet_i_bits_gh_backup(fetch_buffer_io_bpu_inst_packet_i_bits_gh_backup),
    .io_bpu_inst_packet_i_bits_valid_mask_0(fetch_buffer_io_bpu_inst_packet_i_bits_valid_mask_0),
    .io_bpu_inst_packet_i_bits_valid_mask_1(fetch_buffer_io_bpu_inst_packet_i_bits_valid_mask_1),
    .io_bpu_inst_packet_i_bits_valid_mask_2(fetch_buffer_io_bpu_inst_packet_i_bits_valid_mask_2),
    .io_bpu_inst_packet_i_bits_valid_mask_3(fetch_buffer_io_bpu_inst_packet_i_bits_valid_mask_3),
    .io_bpu_inst_packet_i_bits_valid_mask_4(fetch_buffer_io_bpu_inst_packet_i_bits_valid_mask_4),
    .io_bpu_inst_packet_i_bits_valid_mask_5(fetch_buffer_io_bpu_inst_packet_i_bits_valid_mask_5),
    .io_bpu_inst_packet_i_bits_valid_mask_6(fetch_buffer_io_bpu_inst_packet_i_bits_valid_mask_6),
    .io_bpu_inst_packet_i_bits_valid_mask_7(fetch_buffer_io_bpu_inst_packet_i_bits_valid_mask_7),
    .io_bpu_inst_packet_i_bits_predict_mask_0(fetch_buffer_io_bpu_inst_packet_i_bits_predict_mask_0),
    .io_bpu_inst_packet_i_bits_predict_mask_1(fetch_buffer_io_bpu_inst_packet_i_bits_predict_mask_1),
    .io_bpu_inst_packet_i_bits_predict_mask_2(fetch_buffer_io_bpu_inst_packet_i_bits_predict_mask_2),
    .io_bpu_inst_packet_i_bits_predict_mask_3(fetch_buffer_io_bpu_inst_packet_i_bits_predict_mask_3),
    .io_bpu_inst_packet_i_bits_predict_mask_4(fetch_buffer_io_bpu_inst_packet_i_bits_predict_mask_4),
    .io_bpu_inst_packet_i_bits_predict_mask_5(fetch_buffer_io_bpu_inst_packet_i_bits_predict_mask_5),
    .io_bpu_inst_packet_i_bits_predict_mask_6(fetch_buffer_io_bpu_inst_packet_i_bits_predict_mask_6),
    .io_bpu_inst_packet_i_bits_predict_mask_7(fetch_buffer_io_bpu_inst_packet_i_bits_predict_mask_7),
    .io_inst_bank_valid(fetch_buffer_io_inst_bank_valid),
    .io_inst_bank_bits_data_0_inst(fetch_buffer_io_inst_bank_bits_data_0_inst),
    .io_inst_bank_bits_data_0_inst_addr(fetch_buffer_io_inst_bank_bits_data_0_inst_addr),
    .io_inst_bank_bits_data_0_gh_backup(fetch_buffer_io_inst_bank_bits_data_0_gh_backup),
    .io_inst_bank_bits_data_0_is_valid(fetch_buffer_io_inst_bank_bits_data_0_is_valid),
    .io_inst_bank_bits_data_0_predict_taken(fetch_buffer_io_inst_bank_bits_data_0_predict_taken),
    .io_inst_bank_bits_data_1_inst(fetch_buffer_io_inst_bank_bits_data_1_inst),
    .io_inst_bank_bits_data_1_inst_addr(fetch_buffer_io_inst_bank_bits_data_1_inst_addr),
    .io_inst_bank_bits_data_1_gh_backup(fetch_buffer_io_inst_bank_bits_data_1_gh_backup),
    .io_inst_bank_bits_data_1_is_valid(fetch_buffer_io_inst_bank_bits_data_1_is_valid),
    .io_inst_bank_bits_data_1_predict_taken(fetch_buffer_io_inst_bank_bits_data_1_predict_taken),
    .io_fb_resp_deq_valid_0(fetch_buffer_io_fb_resp_deq_valid_0),
    .io_fb_resp_deq_valid_1(fetch_buffer_io_fb_resp_deq_valid_1),
    .io_clear_i(fetch_buffer_io_clear_i)
  );
  assign io_fb_inst_bank_o_valid = fetch_buffer_io_inst_bank_valid; // @[Ifu.scala 62:21]
  assign io_fb_inst_bank_o_bits_data_0_inst = fetch_buffer_io_inst_bank_bits_data_0_inst; // @[Ifu.scala 62:21]
  assign io_fb_inst_bank_o_bits_data_0_inst_addr = fetch_buffer_io_inst_bank_bits_data_0_inst_addr; // @[Ifu.scala 62:21]
  assign io_fb_inst_bank_o_bits_data_0_gh_backup = fetch_buffer_io_inst_bank_bits_data_0_gh_backup; // @[Ifu.scala 62:21]
  assign io_fb_inst_bank_o_bits_data_0_is_valid = fetch_buffer_io_inst_bank_bits_data_0_is_valid; // @[Ifu.scala 62:21]
  assign io_fb_inst_bank_o_bits_data_0_predict_taken = fetch_buffer_io_inst_bank_bits_data_0_predict_taken; // @[Ifu.scala 62:21]
  assign io_fb_inst_bank_o_bits_data_1_inst = fetch_buffer_io_inst_bank_bits_data_1_inst; // @[Ifu.scala 62:21]
  assign io_fb_inst_bank_o_bits_data_1_inst_addr = fetch_buffer_io_inst_bank_bits_data_1_inst_addr; // @[Ifu.scala 62:21]
  assign io_fb_inst_bank_o_bits_data_1_gh_backup = fetch_buffer_io_inst_bank_bits_data_1_gh_backup; // @[Ifu.scala 62:21]
  assign io_fb_inst_bank_o_bits_data_1_is_valid = fetch_buffer_io_inst_bank_bits_data_1_is_valid; // @[Ifu.scala 62:21]
  assign io_fb_inst_bank_o_bits_data_1_predict_taken = fetch_buffer_io_inst_bank_bits_data_1_predict_taken; // @[Ifu.scala 62:21]
  assign io_icache_io_read_req_valid = icache_io_io_read_req_valid; // @[Ifu.scala 53:24]
  assign io_icache_io_read_req_bits_addr = icache_io_io_read_req_bits_addr; // @[Ifu.scala 53:24]
  assign io_icache_debug_state = icache_io_icache_debug_state; // @[Ifu.scala 65:18]
  assign io_icache_debug_hit_cache = icache_io_icache_debug_hit_cache; // @[Ifu.scala 65:18]
  assign io_icache_debug_cache_we = icache_io_icache_debug_cache_we; // @[Ifu.scala 65:18]
  assign io_icache_debug_cache_read_tag = icache_io_icache_debug_cache_read_tag; // @[Ifu.scala 65:18]
  assign io_icache_debug_icache_req_valid = icache_io_icache_debug_icache_req_valid; // @[Ifu.scala 65:18]
  assign io_icache_debug_icache_req_bits_addr = icache_io_icache_debug_icache_req_bits_addr; // @[Ifu.scala 65:18]
  assign io_bpu_debug_branch_mask = bpu_io_bpu_debug_branch_mask; // @[Ifu.scala 66:15]
  assign io_bpu_debug_fetched_mask = bpu_io_bpu_debug_fetched_mask; // @[Ifu.scala 66:15]
  assign io_bpu_debug_predict_branch = bpu_io_bpu_debug_predict_branch; // @[Ifu.scala 66:15]
  assign io_bpu_debug_predict_addr = bpu_io_bpu_debug_predict_addr; // @[Ifu.scala 66:15]
  assign io_bpu_debug_is_taken = bpu_io_bpu_debug_is_taken; // @[Ifu.scala 66:15]
  assign io_bpu_debug_take_delay = bpu_io_bpu_debug_take_delay; // @[Ifu.scala 66:15]
  assign io_bpu_debug_inst_packet_0 = bpu_io_bpu_debug_inst_packet_0; // @[Ifu.scala 66:15]
  assign io_bpu_debug_inst_packet_1 = bpu_io_bpu_debug_inst_packet_1; // @[Ifu.scala 66:15]
  assign io_bpu_debug_inst_packet_2 = bpu_io_bpu_debug_inst_packet_2; // @[Ifu.scala 66:15]
  assign io_bpu_debug_inst_packet_3 = bpu_io_bpu_debug_inst_packet_3; // @[Ifu.scala 66:15]
  assign io_bpu_debug_inst_packet_4 = bpu_io_bpu_debug_inst_packet_4; // @[Ifu.scala 66:15]
  assign io_bpu_debug_inst_packet_5 = bpu_io_bpu_debug_inst_packet_5; // @[Ifu.scala 66:15]
  assign io_bpu_debug_inst_packet_6 = bpu_io_bpu_debug_inst_packet_6; // @[Ifu.scala 66:15]
  assign io_bpu_debug_inst_packet_7 = bpu_io_bpu_debug_inst_packet_7; // @[Ifu.scala 66:15]
  assign bpu_clock = clock;
  assign bpu_reset = reset;
  assign bpu_io_inst_packet_i_valid = icache_io_icache_resp_valid; // @[Ifu.scala 52:25]
  assign bpu_io_inst_packet_i_bits_data_0 = icache_io_icache_resp_bits_data_0; // @[Ifu.scala 52:25]
  assign bpu_io_inst_packet_i_bits_data_1 = icache_io_icache_resp_bits_data_1; // @[Ifu.scala 52:25]
  assign bpu_io_inst_packet_i_bits_data_2 = icache_io_icache_resp_bits_data_2; // @[Ifu.scala 52:25]
  assign bpu_io_inst_packet_i_bits_data_3 = icache_io_icache_resp_bits_data_3; // @[Ifu.scala 52:25]
  assign bpu_io_inst_packet_i_bits_data_4 = icache_io_icache_resp_bits_data_4; // @[Ifu.scala 52:25]
  assign bpu_io_inst_packet_i_bits_data_5 = icache_io_icache_resp_bits_data_5; // @[Ifu.scala 52:25]
  assign bpu_io_inst_packet_i_bits_data_6 = icache_io_icache_resp_bits_data_6; // @[Ifu.scala 52:25]
  assign bpu_io_inst_packet_i_bits_data_7 = icache_io_icache_resp_bits_data_7; // @[Ifu.scala 52:25]
  assign bpu_io_inst_packet_i_bits_addr = icache_io_icache_resp_bits_addr; // @[Ifu.scala 52:25]
  assign bpu_io_bpu_inst_packet_o_ready = fetch_buffer_io_bpu_inst_packet_i_ready; // @[Ifu.scala 57:28]
  assign bpu_io_branch_info_i_valid = io_ex_branch_info_i_valid; // @[Ifu.scala 58:24]
  assign bpu_io_branch_info_i_bits_inst_addr = io_ex_branch_info_i_bits_inst_addr; // @[Ifu.scala 58:24]
  assign bpu_io_branch_info_i_bits_gh_update = io_ex_branch_info_i_bits_gh_update; // @[Ifu.scala 58:24]
  assign bpu_io_branch_info_i_bits_is_branch = io_ex_branch_info_i_bits_is_branch; // @[Ifu.scala 58:24]
  assign bpu_io_branch_info_i_bits_is_taken = io_ex_branch_info_i_bits_is_taken; // @[Ifu.scala 58:24]
  assign bpu_io_branch_info_i_bits_predict_miss = io_ex_branch_info_i_bits_predict_miss; // @[Ifu.scala 58:24]
  assign bpu_io_is_delay = taking_delay; // @[Ifu.scala 56:18]
  assign bpu_io_need_flush = io_ex_branch_info_i_valid & io_ex_branch_info_i_bits_predict_miss; // @[Ifu.scala 26:44]
  assign icache_clock = clock;
  assign icache_reset = reset;
  assign icache_io_icache_req_valid = ~redirect; // @[Ifu.scala 51:33]
  assign icache_io_icache_req_bits_addr = pc; // @[Ifu.scala 50:34]
  assign icache_io_io_read_req_ready = io_icache_io_read_req_ready; // @[Ifu.scala 53:24]
  assign icache_io_io_read_resp_bits_data = io_icache_io_read_resp_bits_data; // @[Ifu.scala 54:25]
  assign fetch_buffer_clock = clock;
  assign fetch_buffer_reset = reset;
  assign fetch_buffer_io_bpu_inst_packet_i_valid = bpu_io_bpu_inst_packet_o_valid; // @[Ifu.scala 57:28]
  assign fetch_buffer_io_bpu_inst_packet_i_bits_data_0 = bpu_io_bpu_inst_packet_o_bits_data_0; // @[Ifu.scala 57:28]
  assign fetch_buffer_io_bpu_inst_packet_i_bits_data_1 = bpu_io_bpu_inst_packet_o_bits_data_1; // @[Ifu.scala 57:28]
  assign fetch_buffer_io_bpu_inst_packet_i_bits_data_2 = bpu_io_bpu_inst_packet_o_bits_data_2; // @[Ifu.scala 57:28]
  assign fetch_buffer_io_bpu_inst_packet_i_bits_data_3 = bpu_io_bpu_inst_packet_o_bits_data_3; // @[Ifu.scala 57:28]
  assign fetch_buffer_io_bpu_inst_packet_i_bits_data_4 = bpu_io_bpu_inst_packet_o_bits_data_4; // @[Ifu.scala 57:28]
  assign fetch_buffer_io_bpu_inst_packet_i_bits_data_5 = bpu_io_bpu_inst_packet_o_bits_data_5; // @[Ifu.scala 57:28]
  assign fetch_buffer_io_bpu_inst_packet_i_bits_data_6 = bpu_io_bpu_inst_packet_o_bits_data_6; // @[Ifu.scala 57:28]
  assign fetch_buffer_io_bpu_inst_packet_i_bits_data_7 = bpu_io_bpu_inst_packet_o_bits_data_7; // @[Ifu.scala 57:28]
  assign fetch_buffer_io_bpu_inst_packet_i_bits_addr = bpu_io_bpu_inst_packet_o_bits_addr; // @[Ifu.scala 57:28]
  assign fetch_buffer_io_bpu_inst_packet_i_bits_gh_backup = bpu_io_bpu_inst_packet_o_bits_gh_backup; // @[Ifu.scala 57:28]
  assign fetch_buffer_io_bpu_inst_packet_i_bits_valid_mask_0 = bpu_io_bpu_inst_packet_o_bits_valid_mask_0; // @[Ifu.scala 57:28]
  assign fetch_buffer_io_bpu_inst_packet_i_bits_valid_mask_1 = bpu_io_bpu_inst_packet_o_bits_valid_mask_1; // @[Ifu.scala 57:28]
  assign fetch_buffer_io_bpu_inst_packet_i_bits_valid_mask_2 = bpu_io_bpu_inst_packet_o_bits_valid_mask_2; // @[Ifu.scala 57:28]
  assign fetch_buffer_io_bpu_inst_packet_i_bits_valid_mask_3 = bpu_io_bpu_inst_packet_o_bits_valid_mask_3; // @[Ifu.scala 57:28]
  assign fetch_buffer_io_bpu_inst_packet_i_bits_valid_mask_4 = bpu_io_bpu_inst_packet_o_bits_valid_mask_4; // @[Ifu.scala 57:28]
  assign fetch_buffer_io_bpu_inst_packet_i_bits_valid_mask_5 = bpu_io_bpu_inst_packet_o_bits_valid_mask_5; // @[Ifu.scala 57:28]
  assign fetch_buffer_io_bpu_inst_packet_i_bits_valid_mask_6 = bpu_io_bpu_inst_packet_o_bits_valid_mask_6; // @[Ifu.scala 57:28]
  assign fetch_buffer_io_bpu_inst_packet_i_bits_valid_mask_7 = bpu_io_bpu_inst_packet_o_bits_valid_mask_7; // @[Ifu.scala 57:28]
  assign fetch_buffer_io_bpu_inst_packet_i_bits_predict_mask_0 = bpu_io_bpu_inst_packet_o_bits_predict_mask_0; // @[Ifu.scala 57:28]
  assign fetch_buffer_io_bpu_inst_packet_i_bits_predict_mask_1 = bpu_io_bpu_inst_packet_o_bits_predict_mask_1; // @[Ifu.scala 57:28]
  assign fetch_buffer_io_bpu_inst_packet_i_bits_predict_mask_2 = bpu_io_bpu_inst_packet_o_bits_predict_mask_2; // @[Ifu.scala 57:28]
  assign fetch_buffer_io_bpu_inst_packet_i_bits_predict_mask_3 = bpu_io_bpu_inst_packet_o_bits_predict_mask_3; // @[Ifu.scala 57:28]
  assign fetch_buffer_io_bpu_inst_packet_i_bits_predict_mask_4 = bpu_io_bpu_inst_packet_o_bits_predict_mask_4; // @[Ifu.scala 57:28]
  assign fetch_buffer_io_bpu_inst_packet_i_bits_predict_mask_5 = bpu_io_bpu_inst_packet_o_bits_predict_mask_5; // @[Ifu.scala 57:28]
  assign fetch_buffer_io_bpu_inst_packet_i_bits_predict_mask_6 = bpu_io_bpu_inst_packet_o_bits_predict_mask_6; // @[Ifu.scala 57:28]
  assign fetch_buffer_io_bpu_inst_packet_i_bits_predict_mask_7 = bpu_io_bpu_inst_packet_o_bits_predict_mask_7; // @[Ifu.scala 57:28]
  assign fetch_buffer_io_fb_resp_deq_valid_0 = io_fb_resp_deq_valid_0; // @[Ifu.scala 63:13]
  assign fetch_buffer_io_fb_resp_deq_valid_1 = io_fb_resp_deq_valid_1; // @[Ifu.scala 63:13]
  assign fetch_buffer_io_clear_i = io_ex_branch_info_i_valid & io_ex_branch_info_i_bits_predict_miss; // @[Ifu.scala 26:44]
  always @(posedge clock) begin
    if (reset) begin // @[Ifu.scala 23:30]
      pc <= 32'h80000000; // @[Ifu.scala 23:30]
    end else if (redirect) begin // @[Ifu.scala 31:18]
      pc <= io_ex_branch_info_i_bits_target_addr; // @[Ifu.scala 32:8]
    end else if (!(stop_fetch)) begin // @[Ifu.scala 34:25]
      if (taking_delay) begin // @[Ifu.scala 36:28]
        pc <= delay_target_addr; // @[Ifu.scala 37:8]
      end else begin
        pc <= _GEN_1;
      end
    end
    if (reset) begin // @[Ifu.scala 28:34]
      taking_delay <= 1'h0; // @[Ifu.scala 28:34]
    end else if (redirect) begin // @[Ifu.scala 31:18]
      taking_delay <= 1'h0; // @[Ifu.scala 33:18]
    end else if (!(stop_fetch)) begin // @[Ifu.scala 34:25]
      if (taking_delay) begin // @[Ifu.scala 36:28]
        taking_delay <= 1'h0; // @[Ifu.scala 38:18]
      end else begin
        taking_delay <= _GEN_2;
      end
    end
    if (reset) begin // @[Ifu.scala 29:34]
      delay_target_addr <= 32'h0; // @[Ifu.scala 29:34]
    end else if (!(redirect)) begin // @[Ifu.scala 31:18]
      if (!(stop_fetch)) begin // @[Ifu.scala 34:25]
        if (!(taking_delay)) begin // @[Ifu.scala 36:28]
          delay_target_addr <= _GEN_3;
        end
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  pc = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  taking_delay = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  delay_target_addr = _RAND_2[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Decode(
  input         clock,
  input         reset,
  input         io_fb_inst_bank_valid,
  input  [31:0] io_fb_inst_bank_bits_data_0_inst,
  input  [31:0] io_fb_inst_bank_bits_data_0_inst_addr,
  input  [3:0]  io_fb_inst_bank_bits_data_0_gh_backup,
  input         io_fb_inst_bank_bits_data_0_is_valid,
  input         io_fb_inst_bank_bits_data_0_predict_taken,
  input  [31:0] io_fb_inst_bank_bits_data_1_inst,
  input  [31:0] io_fb_inst_bank_bits_data_1_inst_addr,
  input  [3:0]  io_fb_inst_bank_bits_data_1_gh_backup,
  input         io_fb_inst_bank_bits_data_1_is_valid,
  input         io_fb_inst_bank_bits_data_1_predict_taken,
  output        io_fb_resp_deq_valid_0,
  output        io_fb_resp_deq_valid_1,
  output        io_rob_allocate_allocate_req_valid,
  output        io_rob_allocate_allocate_req_bits_0,
  output        io_rob_allocate_allocate_req_bits_1,
  output        io_rob_allocate_allocate_info_valid,
  output [2:0]  io_rob_allocate_allocate_info_bits_0_rob_idx,
  output        io_rob_allocate_allocate_info_bits_0_inst_valid,
  output [31:0] io_rob_allocate_allocate_info_bits_0_inst_addr,
  output [5:0]  io_rob_allocate_allocate_info_bits_0_uop,
  output [2:0]  io_rob_allocate_allocate_info_bits_0_unit_sel,
  output        io_rob_allocate_allocate_info_bits_0_need_imm,
  output [31:0] io_rob_allocate_allocate_info_bits_0_commit_addr,
  output [3:0]  io_rob_allocate_allocate_info_bits_0_gh_info,
  output [31:0] io_rob_allocate_allocate_info_bits_0_imm_data,
  output        io_rob_allocate_allocate_info_bits_0_flush_on_commit,
  output        io_rob_allocate_allocate_info_bits_0_predict_taken,
  output [2:0]  io_rob_allocate_allocate_info_bits_1_rob_idx,
  output        io_rob_allocate_allocate_info_bits_1_inst_valid,
  output [31:0] io_rob_allocate_allocate_info_bits_1_inst_addr,
  output [5:0]  io_rob_allocate_allocate_info_bits_1_uop,
  output [2:0]  io_rob_allocate_allocate_info_bits_1_unit_sel,
  output        io_rob_allocate_allocate_info_bits_1_need_imm,
  output [31:0] io_rob_allocate_allocate_info_bits_1_commit_addr,
  output [3:0]  io_rob_allocate_allocate_info_bits_1_gh_info,
  output [31:0] io_rob_allocate_allocate_info_bits_1_imm_data,
  output        io_rob_allocate_allocate_info_bits_1_flush_on_commit,
  output        io_rob_allocate_allocate_info_bits_1_predict_taken,
  input         io_rob_allocate_allocate_resp_valid,
  input  [2:0]  io_rob_allocate_allocate_resp_bits_rob_idx_0,
  input  [2:0]  io_rob_allocate_allocate_resp_bits_rob_idx_1,
  input         io_rob_allocate_allocate_resp_bits_enq_valid_mask_0,
  input         io_rob_allocate_allocate_resp_bits_enq_valid_mask_1,
  output        io_rename_info_valid,
  output        io_rename_info_bits_0_is_valid,
  output [4:0]  io_rename_info_bits_0_op1_addr,
  output [4:0]  io_rename_info_bits_0_op2_addr,
  output [4:0]  io_rename_info_bits_0_des_addr,
  output [2:0]  io_rename_info_bits_0_des_rob,
  output        io_rename_info_bits_1_is_valid,
  output [4:0]  io_rename_info_bits_1_op1_addr,
  output [4:0]  io_rename_info_bits_1_op2_addr,
  output [4:0]  io_rename_info_bits_1_des_addr,
  output [2:0]  io_rename_info_bits_1_des_rob,
  input         io_need_flush
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
`endif // RANDOMIZE_REG_INIT
  wire [31:0] _decoder_T = io_fb_inst_bank_bits_data_0_inst & 32'hfc0007ff; // @[Lookup.scala 31:38]
  wire  _decoder_T_1 = 32'h20 == _decoder_T; // @[Lookup.scala 31:38]
  wire [31:0] _decoder_T_2 = io_fb_inst_bank_bits_data_0_inst & 32'hfc000000; // @[Lookup.scala 31:38]
  wire  _decoder_T_3 = 32'h20000000 == _decoder_T_2; // @[Lookup.scala 31:38]
  wire  _decoder_T_5 = 32'h21 == _decoder_T; // @[Lookup.scala 31:38]
  wire  _decoder_T_7 = 32'h24000000 == _decoder_T_2; // @[Lookup.scala 31:38]
  wire  _decoder_T_9 = 32'h22 == _decoder_T; // @[Lookup.scala 31:38]
  wire  _decoder_T_11 = 32'h23 == _decoder_T; // @[Lookup.scala 31:38]
  wire  _decoder_T_13 = 32'h2a == _decoder_T; // @[Lookup.scala 31:38]
  wire  _decoder_T_15 = 32'h28000000 == _decoder_T_2; // @[Lookup.scala 31:38]
  wire  _decoder_T_17 = 32'h2b == _decoder_T; // @[Lookup.scala 31:38]
  wire  _decoder_T_19 = 32'h2c000000 == _decoder_T_2; // @[Lookup.scala 31:38]
  wire  _decoder_T_21 = 32'h70000002 == _decoder_T; // @[Lookup.scala 31:38]
  wire [31:0] _decoder_T_22 = io_fb_inst_bank_bits_data_0_inst & 32'hfc00ffff; // @[Lookup.scala 31:38]
  wire  _decoder_T_23 = 32'h1a == _decoder_T_22; // @[Lookup.scala 31:38]
  wire  _decoder_T_25 = 32'h1b == _decoder_T_22; // @[Lookup.scala 31:38]
  wire  _decoder_T_27 = 32'h18 == _decoder_T_22; // @[Lookup.scala 31:38]
  wire  _decoder_T_29 = 32'h19 == _decoder_T_22; // @[Lookup.scala 31:38]
  wire [31:0] _decoder_T_30 = io_fb_inst_bank_bits_data_0_inst & 32'hffff07ff; // @[Lookup.scala 31:38]
  wire  _decoder_T_31 = 32'h10 == _decoder_T_30; // @[Lookup.scala 31:38]
  wire  _decoder_T_33 = 32'h12 == _decoder_T_30; // @[Lookup.scala 31:38]
  wire [31:0] _decoder_T_34 = io_fb_inst_bank_bits_data_0_inst & 32'hfc1fffff; // @[Lookup.scala 31:38]
  wire  _decoder_T_35 = 32'h11 == _decoder_T_34; // @[Lookup.scala 31:38]
  wire  _decoder_T_37 = 32'h13 == _decoder_T_34; // @[Lookup.scala 31:38]
  wire  _decoder_T_39 = 32'h24 == _decoder_T; // @[Lookup.scala 31:38]
  wire  _decoder_T_41 = 32'h30000000 == _decoder_T_2; // @[Lookup.scala 31:38]
  wire [31:0] _decoder_T_42 = io_fb_inst_bank_bits_data_0_inst & 32'hffe00000; // @[Lookup.scala 31:38]
  wire  _decoder_T_43 = 32'h3c000000 == _decoder_T_42; // @[Lookup.scala 31:38]
  wire  _decoder_T_45 = 32'h27 == _decoder_T; // @[Lookup.scala 31:38]
  wire  _decoder_T_47 = 32'h25 == _decoder_T; // @[Lookup.scala 31:38]
  wire  _decoder_T_49 = 32'h34000000 == _decoder_T_2; // @[Lookup.scala 31:38]
  wire  _decoder_T_51 = 32'h26 == _decoder_T; // @[Lookup.scala 31:38]
  wire  _decoder_T_53 = 32'h38000000 == _decoder_T_2; // @[Lookup.scala 31:38]
  wire  _decoder_T_55 = 32'h4 == _decoder_T; // @[Lookup.scala 31:38]
  wire [31:0] _decoder_T_56 = io_fb_inst_bank_bits_data_0_inst & 32'hffe0003f; // @[Lookup.scala 31:38]
  wire  _decoder_T_57 = 32'h0 == _decoder_T_56; // @[Lookup.scala 31:38]
  wire  _decoder_T_59 = 32'h7 == _decoder_T; // @[Lookup.scala 31:38]
  wire  _decoder_T_61 = 32'h3 == _decoder_T_56; // @[Lookup.scala 31:38]
  wire  _decoder_T_63 = 32'h6 == _decoder_T; // @[Lookup.scala 31:38]
  wire  _decoder_T_65 = 32'h2 == _decoder_T_56; // @[Lookup.scala 31:38]
  wire  _decoder_T_67 = 32'h10000000 == _decoder_T_2; // @[Lookup.scala 31:38]
  wire  _decoder_T_69 = 32'h14000000 == _decoder_T_2; // @[Lookup.scala 31:38]
  wire [31:0] _decoder_T_70 = io_fb_inst_bank_bits_data_0_inst & 32'hfc1f0000; // @[Lookup.scala 31:38]
  wire  _decoder_T_71 = 32'h4010000 == _decoder_T_70; // @[Lookup.scala 31:38]
  wire  _decoder_T_73 = 32'h1c000000 == _decoder_T_70; // @[Lookup.scala 31:38]
  wire  _decoder_T_75 = 32'h18000000 == _decoder_T_70; // @[Lookup.scala 31:38]
  wire  _decoder_T_77 = 32'h4000000 == _decoder_T_70; // @[Lookup.scala 31:38]
  wire  _decoder_T_83 = 32'h8000000 == _decoder_T_2; // @[Lookup.scala 31:38]
  wire  _decoder_T_85 = 32'hc000000 == _decoder_T_2; // @[Lookup.scala 31:38]
  wire  _decoder_T_87 = 32'h8 == _decoder_T_34; // @[Lookup.scala 31:38]
  wire [31:0] _decoder_T_88 = io_fb_inst_bank_bits_data_0_inst & 32'hfc1f07ff; // @[Lookup.scala 31:38]
  wire  _decoder_T_89 = 32'h9 == _decoder_T_88; // @[Lookup.scala 31:38]
  wire  _decoder_T_91 = 32'hc == io_fb_inst_bank_bits_data_0_inst; // @[Lookup.scala 31:38]
  wire [31:0] _decoder_T_92 = io_fb_inst_bank_bits_data_0_inst & 32'hfc00003f; // @[Lookup.scala 31:38]
  wire  _decoder_T_93 = 32'hd == _decoder_T_92; // @[Lookup.scala 31:38]
  wire  _decoder_T_95 = 32'h42000018 == io_fb_inst_bank_bits_data_0_inst; // @[Lookup.scala 31:38]
  wire [31:0] _decoder_T_96 = io_fb_inst_bank_bits_data_0_inst & 32'hffe007ff; // @[Lookup.scala 31:38]
  wire  _decoder_T_97 = 32'h40000000 == _decoder_T_96; // @[Lookup.scala 31:38]
  wire  _decoder_T_99 = 32'h40800000 == _decoder_T_96; // @[Lookup.scala 31:38]
  wire  _decoder_T_101 = 32'h80000000 == _decoder_T_2; // @[Lookup.scala 31:38]
  wire  _decoder_T_103 = 32'h84000000 == _decoder_T_2; // @[Lookup.scala 31:38]
  wire  _decoder_T_105 = 32'h8c000000 == _decoder_T_2; // @[Lookup.scala 31:38]
  wire  _decoder_T_107 = 32'h90000000 == _decoder_T_2; // @[Lookup.scala 31:38]
  wire  _decoder_T_109 = 32'h94000000 == _decoder_T_2; // @[Lookup.scala 31:38]
  wire  _decoder_T_111 = 32'ha0000000 == _decoder_T_2; // @[Lookup.scala 31:38]
  wire  _decoder_T_113 = 32'ha4000000 == _decoder_T_2; // @[Lookup.scala 31:38]
  wire  _decoder_T_115 = 32'hac000000 == _decoder_T_2; // @[Lookup.scala 31:38]
  wire [5:0] _decoder_T_116 = _decoder_T_115 ? 6'h24 : 6'h0; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_117 = _decoder_T_113 ? 6'h25 : _decoder_T_116; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_118 = _decoder_T_111 ? 6'h26 : _decoder_T_117; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_119 = _decoder_T_109 ? 6'h29 : _decoder_T_118; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_120 = _decoder_T_107 ? 6'h2b : _decoder_T_119; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_121 = _decoder_T_105 ? 6'h27 : _decoder_T_120; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_122 = _decoder_T_103 ? 6'h28 : _decoder_T_121; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_123 = _decoder_T_101 ? 6'h2a : _decoder_T_122; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_124 = _decoder_T_99 ? 6'h2c : _decoder_T_123; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_125 = _decoder_T_97 ? 6'h2d : _decoder_T_124; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_126 = _decoder_T_95 ? 6'h2f : _decoder_T_125; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_127 = _decoder_T_93 ? 6'h30 : _decoder_T_126; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_128 = _decoder_T_91 ? 6'h2e : _decoder_T_127; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_129 = _decoder_T_89 ? 6'h1b : _decoder_T_128; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_130 = _decoder_T_87 ? 6'h1a : _decoder_T_129; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_131 = _decoder_T_85 ? 6'h19 : _decoder_T_130; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_132 = _decoder_T_83 ? 6'h18 : _decoder_T_131; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_133 = _decoder_T_75 ? 6'h23 : _decoder_T_132; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_134 = _decoder_T_71 ? 6'h22 : _decoder_T_133; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_135 = _decoder_T_77 ? 6'h20 : _decoder_T_134; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_136 = _decoder_T_75 ? 6'h1e : _decoder_T_135; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_137 = _decoder_T_73 ? 6'h1f : _decoder_T_136; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_138 = _decoder_T_71 ? 6'h21 : _decoder_T_137; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_139 = _decoder_T_69 ? 6'h1d : _decoder_T_138; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_140 = _decoder_T_67 ? 6'h1c : _decoder_T_139; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_141 = _decoder_T_65 ? 6'h6 : _decoder_T_140; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_142 = _decoder_T_63 ? 6'h6 : _decoder_T_141; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_143 = _decoder_T_61 ? 6'h7 : _decoder_T_142; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_144 = _decoder_T_59 ? 6'h7 : _decoder_T_143; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_145 = _decoder_T_57 ? 6'h5 : _decoder_T_144; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_146 = _decoder_T_55 ? 6'h5 : _decoder_T_145; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_147 = _decoder_T_53 ? 6'ha : _decoder_T_146; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_148 = _decoder_T_51 ? 6'ha : _decoder_T_147; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_149 = _decoder_T_49 ? 6'hb : _decoder_T_148; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_150 = _decoder_T_47 ? 6'hb : _decoder_T_149; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_151 = _decoder_T_45 ? 6'he : _decoder_T_150; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_152 = _decoder_T_43 ? 6'hd : _decoder_T_151; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_153 = _decoder_T_41 ? 6'hc : _decoder_T_152; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_154 = _decoder_T_39 ? 6'hc : _decoder_T_153; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_155 = _decoder_T_37 ? 6'h17 : _decoder_T_154; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_156 = _decoder_T_35 ? 6'h16 : _decoder_T_155; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_157 = _decoder_T_33 ? 6'h15 : _decoder_T_156; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_158 = _decoder_T_31 ? 6'h14 : _decoder_T_157; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_159 = _decoder_T_29 ? 6'h11 : _decoder_T_158; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_160 = _decoder_T_27 ? 6'h10 : _decoder_T_159; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_161 = _decoder_T_25 ? 6'h13 : _decoder_T_160; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_162 = _decoder_T_23 ? 6'h12 : _decoder_T_161; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_163 = _decoder_T_21 ? 6'hf : _decoder_T_162; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_164 = _decoder_T_19 ? 6'h9 : _decoder_T_163; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_165 = _decoder_T_17 ? 6'h9 : _decoder_T_164; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_166 = _decoder_T_15 ? 6'h8 : _decoder_T_165; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_167 = _decoder_T_13 ? 6'h8 : _decoder_T_166; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_168 = _decoder_T_11 ? 6'h4 : _decoder_T_167; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_169 = _decoder_T_9 ? 6'h3 : _decoder_T_168; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_170 = _decoder_T_7 ? 6'h2 : _decoder_T_169; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_171 = _decoder_T_5 ? 6'h2 : _decoder_T_170; // @[Lookup.scala 33:37]
  wire [1:0] _decoder_T_173 = _decoder_T_115 ? 2'h3 : 2'h0; // @[Lookup.scala 33:37]
  wire [1:0] _decoder_T_174 = _decoder_T_113 ? 2'h3 : _decoder_T_173; // @[Lookup.scala 33:37]
  wire [1:0] _decoder_T_175 = _decoder_T_111 ? 2'h3 : _decoder_T_174; // @[Lookup.scala 33:37]
  wire [1:0] _decoder_T_176 = _decoder_T_109 ? 2'h3 : _decoder_T_175; // @[Lookup.scala 33:37]
  wire [1:0] _decoder_T_177 = _decoder_T_107 ? 2'h3 : _decoder_T_176; // @[Lookup.scala 33:37]
  wire [1:0] _decoder_T_178 = _decoder_T_105 ? 2'h3 : _decoder_T_177; // @[Lookup.scala 33:37]
  wire [1:0] _decoder_T_179 = _decoder_T_103 ? 2'h3 : _decoder_T_178; // @[Lookup.scala 33:37]
  wire [1:0] _decoder_T_180 = _decoder_T_101 ? 2'h3 : _decoder_T_179; // @[Lookup.scala 33:37]
  wire [1:0] _decoder_T_181 = _decoder_T_99 ? 2'h2 : _decoder_T_180; // @[Lookup.scala 33:37]
  wire [1:0] _decoder_T_182 = _decoder_T_97 ? 2'h2 : _decoder_T_181; // @[Lookup.scala 33:37]
  wire [1:0] _decoder_T_183 = _decoder_T_95 ? 2'h0 : _decoder_T_182; // @[Lookup.scala 33:37]
  wire [1:0] _decoder_T_184 = _decoder_T_93 ? 2'h0 : _decoder_T_183; // @[Lookup.scala 33:37]
  wire [1:0] _decoder_T_185 = _decoder_T_91 ? 2'h0 : _decoder_T_184; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_186 = _decoder_T_89 ? 3'h5 : {{1'd0}, _decoder_T_185}; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_187 = _decoder_T_87 ? 3'h5 : _decoder_T_186; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_188 = _decoder_T_85 ? 3'h5 : _decoder_T_187; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_189 = _decoder_T_83 ? 3'h5 : _decoder_T_188; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_190 = _decoder_T_75 ? 3'h5 : _decoder_T_189; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_191 = _decoder_T_71 ? 3'h5 : _decoder_T_190; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_192 = _decoder_T_77 ? 3'h5 : _decoder_T_191; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_193 = _decoder_T_75 ? 3'h5 : _decoder_T_192; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_194 = _decoder_T_73 ? 3'h5 : _decoder_T_193; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_195 = _decoder_T_71 ? 3'h5 : _decoder_T_194; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_196 = _decoder_T_69 ? 3'h5 : _decoder_T_195; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_197 = _decoder_T_67 ? 3'h5 : _decoder_T_196; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_198 = _decoder_T_65 ? 3'h1 : _decoder_T_197; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_199 = _decoder_T_63 ? 3'h1 : _decoder_T_198; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_200 = _decoder_T_61 ? 3'h1 : _decoder_T_199; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_201 = _decoder_T_59 ? 3'h1 : _decoder_T_200; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_202 = _decoder_T_57 ? 3'h1 : _decoder_T_201; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_203 = _decoder_T_55 ? 3'h1 : _decoder_T_202; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_204 = _decoder_T_53 ? 3'h1 : _decoder_T_203; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_205 = _decoder_T_51 ? 3'h1 : _decoder_T_204; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_206 = _decoder_T_49 ? 3'h1 : _decoder_T_205; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_207 = _decoder_T_47 ? 3'h1 : _decoder_T_206; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_208 = _decoder_T_45 ? 3'h1 : _decoder_T_207; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_209 = _decoder_T_43 ? 3'h1 : _decoder_T_208; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_210 = _decoder_T_41 ? 3'h1 : _decoder_T_209; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_211 = _decoder_T_39 ? 3'h1 : _decoder_T_210; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_212 = _decoder_T_37 ? 3'h4 : _decoder_T_211; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_213 = _decoder_T_35 ? 3'h4 : _decoder_T_212; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_214 = _decoder_T_33 ? 3'h4 : _decoder_T_213; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_215 = _decoder_T_31 ? 3'h4 : _decoder_T_214; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_216 = _decoder_T_29 ? 3'h4 : _decoder_T_215; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_217 = _decoder_T_27 ? 3'h4 : _decoder_T_216; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_218 = _decoder_T_25 ? 3'h4 : _decoder_T_217; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_219 = _decoder_T_23 ? 3'h4 : _decoder_T_218; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_220 = _decoder_T_21 ? 3'h4 : _decoder_T_219; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_221 = _decoder_T_19 ? 3'h1 : _decoder_T_220; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_222 = _decoder_T_17 ? 3'h1 : _decoder_T_221; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_223 = _decoder_T_15 ? 3'h1 : _decoder_T_222; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_224 = _decoder_T_13 ? 3'h1 : _decoder_T_223; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_225 = _decoder_T_11 ? 3'h1 : _decoder_T_224; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_226 = _decoder_T_9 ? 3'h1 : _decoder_T_225; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_227 = _decoder_T_7 ? 3'h1 : _decoder_T_226; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_228 = _decoder_T_5 ? 3'h1 : _decoder_T_227; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_230 = _decoder_T_115 ? 3'h1 : 3'h4; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_231 = _decoder_T_113 ? 3'h1 : _decoder_T_230; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_232 = _decoder_T_111 ? 3'h1 : _decoder_T_231; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_233 = _decoder_T_109 ? 3'h1 : _decoder_T_232; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_234 = _decoder_T_107 ? 3'h1 : _decoder_T_233; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_235 = _decoder_T_105 ? 3'h1 : _decoder_T_234; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_236 = _decoder_T_103 ? 3'h1 : _decoder_T_235; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_237 = _decoder_T_101 ? 3'h1 : _decoder_T_236; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_238 = _decoder_T_99 ? 3'h0 : _decoder_T_237; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_239 = _decoder_T_97 ? 3'h0 : _decoder_T_238; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_240 = _decoder_T_95 ? 3'h4 : _decoder_T_239; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_241 = _decoder_T_93 ? 3'h4 : _decoder_T_240; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_242 = _decoder_T_91 ? 3'h4 : _decoder_T_241; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_243 = _decoder_T_89 ? 3'h4 : _decoder_T_242; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_244 = _decoder_T_87 ? 3'h4 : _decoder_T_243; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_245 = _decoder_T_85 ? 3'h3 : _decoder_T_244; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_246 = _decoder_T_83 ? 3'h3 : _decoder_T_245; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_247 = _decoder_T_75 ? 3'h1 : _decoder_T_246; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_248 = _decoder_T_71 ? 3'h1 : _decoder_T_247; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_249 = _decoder_T_77 ? 3'h1 : _decoder_T_248; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_250 = _decoder_T_75 ? 3'h1 : _decoder_T_249; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_251 = _decoder_T_73 ? 3'h1 : _decoder_T_250; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_252 = _decoder_T_71 ? 3'h1 : _decoder_T_251; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_253 = _decoder_T_69 ? 3'h1 : _decoder_T_252; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_254 = _decoder_T_67 ? 3'h1 : _decoder_T_253; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_255 = _decoder_T_65 ? 3'h2 : _decoder_T_254; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_256 = _decoder_T_63 ? 3'h4 : _decoder_T_255; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_257 = _decoder_T_61 ? 3'h2 : _decoder_T_256; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_258 = _decoder_T_59 ? 3'h4 : _decoder_T_257; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_259 = _decoder_T_57 ? 3'h2 : _decoder_T_258; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_260 = _decoder_T_55 ? 3'h4 : _decoder_T_259; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_261 = _decoder_T_53 ? 3'h0 : _decoder_T_260; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_262 = _decoder_T_51 ? 3'h4 : _decoder_T_261; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_263 = _decoder_T_49 ? 3'h0 : _decoder_T_262; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_264 = _decoder_T_47 ? 3'h4 : _decoder_T_263; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_265 = _decoder_T_45 ? 3'h4 : _decoder_T_264; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_266 = _decoder_T_43 ? 3'h0 : _decoder_T_265; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_267 = _decoder_T_41 ? 3'h0 : _decoder_T_266; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_268 = _decoder_T_39 ? 3'h4 : _decoder_T_267; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_269 = _decoder_T_37 ? 3'h4 : _decoder_T_268; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_270 = _decoder_T_35 ? 3'h4 : _decoder_T_269; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_271 = _decoder_T_33 ? 3'h4 : _decoder_T_270; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_272 = _decoder_T_31 ? 3'h4 : _decoder_T_271; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_273 = _decoder_T_29 ? 3'h4 : _decoder_T_272; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_274 = _decoder_T_27 ? 3'h4 : _decoder_T_273; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_275 = _decoder_T_25 ? 3'h4 : _decoder_T_274; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_276 = _decoder_T_23 ? 3'h4 : _decoder_T_275; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_277 = _decoder_T_21 ? 3'h4 : _decoder_T_276; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_278 = _decoder_T_19 ? 3'h1 : _decoder_T_277; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_279 = _decoder_T_17 ? 3'h4 : _decoder_T_278; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_280 = _decoder_T_15 ? 3'h1 : _decoder_T_279; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_281 = _decoder_T_13 ? 3'h4 : _decoder_T_280; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_282 = _decoder_T_11 ? 3'h4 : _decoder_T_281; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_283 = _decoder_T_9 ? 3'h4 : _decoder_T_282; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_284 = _decoder_T_7 ? 3'h1 : _decoder_T_283; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_285 = _decoder_T_5 ? 3'h4 : _decoder_T_284; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_286 = _decoder_T_3 ? 3'h1 : _decoder_T_285; // @[Lookup.scala 33:37]
  wire [2:0] decoder_2 = _decoder_T_1 ? 3'h4 : _decoder_T_286; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_287 = _decoder_T_115 ? 3'h0 : 3'h4; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_288 = _decoder_T_113 ? 3'h0 : _decoder_T_287; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_289 = _decoder_T_111 ? 3'h0 : _decoder_T_288; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_290 = _decoder_T_109 ? 3'h0 : _decoder_T_289; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_291 = _decoder_T_107 ? 3'h0 : _decoder_T_290; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_292 = _decoder_T_105 ? 3'h0 : _decoder_T_291; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_293 = _decoder_T_103 ? 3'h0 : _decoder_T_292; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_294 = _decoder_T_101 ? 3'h0 : _decoder_T_293; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_295 = _decoder_T_99 ? 3'h1 : _decoder_T_294; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_296 = _decoder_T_97 ? 3'h2 : _decoder_T_295; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_297 = _decoder_T_95 ? 3'h4 : _decoder_T_296; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_298 = _decoder_T_93 ? 3'h4 : _decoder_T_297; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_299 = _decoder_T_91 ? 3'h4 : _decoder_T_298; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_300 = _decoder_T_89 ? 3'h0 : _decoder_T_299; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_301 = _decoder_T_87 ? 3'h0 : _decoder_T_300; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_302 = _decoder_T_85 ? 3'h4 : _decoder_T_301; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_303 = _decoder_T_83 ? 3'h4 : _decoder_T_302; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_304 = _decoder_T_75 ? 3'h0 : _decoder_T_303; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_305 = _decoder_T_71 ? 3'h0 : _decoder_T_304; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_306 = _decoder_T_77 ? 3'h0 : _decoder_T_305; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_307 = _decoder_T_75 ? 3'h0 : _decoder_T_306; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_308 = _decoder_T_73 ? 3'h0 : _decoder_T_307; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_309 = _decoder_T_71 ? 3'h0 : _decoder_T_308; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_310 = _decoder_T_69 ? 3'h0 : _decoder_T_309; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_311 = _decoder_T_67 ? 3'h0 : _decoder_T_310; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_312 = _decoder_T_65 ? 3'h1 : _decoder_T_311; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_313 = _decoder_T_63 ? 3'h1 : _decoder_T_312; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_314 = _decoder_T_61 ? 3'h1 : _decoder_T_313; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_315 = _decoder_T_59 ? 3'h1 : _decoder_T_314; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_316 = _decoder_T_57 ? 3'h1 : _decoder_T_315; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_317 = _decoder_T_55 ? 3'h1 : _decoder_T_316; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_318 = _decoder_T_53 ? 3'h0 : _decoder_T_317; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_319 = _decoder_T_51 ? 3'h0 : _decoder_T_318; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_320 = _decoder_T_49 ? 3'h0 : _decoder_T_319; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_321 = _decoder_T_47 ? 3'h0 : _decoder_T_320; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_322 = _decoder_T_45 ? 3'h0 : _decoder_T_321; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_323 = _decoder_T_43 ? 3'h4 : _decoder_T_322; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_324 = _decoder_T_41 ? 3'h0 : _decoder_T_323; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_325 = _decoder_T_39 ? 3'h0 : _decoder_T_324; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_326 = _decoder_T_37 ? 3'h0 : _decoder_T_325; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_327 = _decoder_T_35 ? 3'h0 : _decoder_T_326; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_328 = _decoder_T_33 ? 3'h4 : _decoder_T_327; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_329 = _decoder_T_31 ? 3'h4 : _decoder_T_328; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_330 = _decoder_T_29 ? 3'h0 : _decoder_T_329; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_331 = _decoder_T_27 ? 3'h0 : _decoder_T_330; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_332 = _decoder_T_25 ? 3'h0 : _decoder_T_331; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_333 = _decoder_T_23 ? 3'h0 : _decoder_T_332; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_334 = _decoder_T_21 ? 3'h0 : _decoder_T_333; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_335 = _decoder_T_19 ? 3'h0 : _decoder_T_334; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_336 = _decoder_T_17 ? 3'h0 : _decoder_T_335; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_337 = _decoder_T_15 ? 3'h0 : _decoder_T_336; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_338 = _decoder_T_13 ? 3'h0 : _decoder_T_337; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_339 = _decoder_T_11 ? 3'h0 : _decoder_T_338; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_340 = _decoder_T_9 ? 3'h0 : _decoder_T_339; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_341 = _decoder_T_7 ? 3'h0 : _decoder_T_340; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_342 = _decoder_T_5 ? 3'h0 : _decoder_T_341; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_343 = _decoder_T_3 ? 3'h0 : _decoder_T_342; // @[Lookup.scala 33:37]
  wire [2:0] decoder_3 = _decoder_T_1 ? 3'h0 : _decoder_T_343; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_347 = _decoder_T_109 ? 3'h4 : _decoder_T_232; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_348 = _decoder_T_107 ? 3'h4 : _decoder_T_347; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_349 = _decoder_T_105 ? 3'h4 : _decoder_T_348; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_350 = _decoder_T_103 ? 3'h4 : _decoder_T_349; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_351 = _decoder_T_101 ? 3'h4 : _decoder_T_350; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_352 = _decoder_T_99 ? 3'h2 : _decoder_T_351; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_353 = _decoder_T_97 ? 3'h4 : _decoder_T_352; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_354 = _decoder_T_95 ? 3'h4 : _decoder_T_353; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_355 = _decoder_T_93 ? 3'h4 : _decoder_T_354; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_356 = _decoder_T_91 ? 3'h4 : _decoder_T_355; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_357 = _decoder_T_89 ? 3'h4 : _decoder_T_356; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_358 = _decoder_T_87 ? 3'h4 : _decoder_T_357; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_359 = _decoder_T_85 ? 3'h4 : _decoder_T_358; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_360 = _decoder_T_83 ? 3'h4 : _decoder_T_359; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_361 = _decoder_T_75 ? 3'h4 : _decoder_T_360; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_362 = _decoder_T_71 ? 3'h4 : _decoder_T_361; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_363 = _decoder_T_77 ? 3'h4 : _decoder_T_362; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_364 = _decoder_T_75 ? 3'h4 : _decoder_T_363; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_365 = _decoder_T_73 ? 3'h4 : _decoder_T_364; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_366 = _decoder_T_71 ? 3'h4 : _decoder_T_365; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_367 = _decoder_T_69 ? 3'h1 : _decoder_T_366; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_368 = _decoder_T_67 ? 3'h1 : _decoder_T_367; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_369 = _decoder_T_65 ? 3'h4 : _decoder_T_368; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_370 = _decoder_T_63 ? 3'h0 : _decoder_T_369; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_371 = _decoder_T_61 ? 3'h4 : _decoder_T_370; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_372 = _decoder_T_59 ? 3'h0 : _decoder_T_371; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_373 = _decoder_T_57 ? 3'h4 : _decoder_T_372; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_374 = _decoder_T_55 ? 3'h0 : _decoder_T_373; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_375 = _decoder_T_53 ? 3'h4 : _decoder_T_374; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_376 = _decoder_T_51 ? 3'h1 : _decoder_T_375; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_377 = _decoder_T_49 ? 3'h4 : _decoder_T_376; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_378 = _decoder_T_47 ? 3'h1 : _decoder_T_377; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_379 = _decoder_T_45 ? 3'h1 : _decoder_T_378; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_380 = _decoder_T_43 ? 3'h4 : _decoder_T_379; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_381 = _decoder_T_41 ? 3'h4 : _decoder_T_380; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_382 = _decoder_T_39 ? 3'h1 : _decoder_T_381; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_383 = _decoder_T_37 ? 3'h4 : _decoder_T_382; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_384 = _decoder_T_35 ? 3'h4 : _decoder_T_383; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_385 = _decoder_T_33 ? 3'h4 : _decoder_T_384; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_386 = _decoder_T_31 ? 3'h4 : _decoder_T_385; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_387 = _decoder_T_29 ? 3'h1 : _decoder_T_386; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_388 = _decoder_T_27 ? 3'h1 : _decoder_T_387; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_389 = _decoder_T_25 ? 3'h1 : _decoder_T_388; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_390 = _decoder_T_23 ? 3'h1 : _decoder_T_389; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_391 = _decoder_T_21 ? 3'h1 : _decoder_T_390; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_392 = _decoder_T_19 ? 3'h4 : _decoder_T_391; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_393 = _decoder_T_17 ? 3'h1 : _decoder_T_392; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_394 = _decoder_T_15 ? 3'h4 : _decoder_T_393; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_395 = _decoder_T_13 ? 3'h1 : _decoder_T_394; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_396 = _decoder_T_11 ? 3'h1 : _decoder_T_395; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_397 = _decoder_T_9 ? 3'h1 : _decoder_T_396; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_398 = _decoder_T_7 ? 3'h4 : _decoder_T_397; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_399 = _decoder_T_5 ? 3'h1 : _decoder_T_398; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_400 = _decoder_T_3 ? 3'h4 : _decoder_T_399; // @[Lookup.scala 33:37]
  wire [2:0] decoder_4 = _decoder_T_1 ? 3'h1 : _decoder_T_400; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_404 = _decoder_T_109 ? 3'h1 : 3'h4; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_405 = _decoder_T_107 ? 3'h1 : _decoder_T_404; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_406 = _decoder_T_105 ? 3'h1 : _decoder_T_405; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_407 = _decoder_T_103 ? 3'h1 : _decoder_T_406; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_408 = _decoder_T_101 ? 3'h1 : _decoder_T_407; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_409 = _decoder_T_99 ? 3'h4 : _decoder_T_408; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_410 = _decoder_T_97 ? 3'h1 : _decoder_T_409; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_411 = _decoder_T_95 ? 3'h4 : _decoder_T_410; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_412 = _decoder_T_93 ? 3'h4 : _decoder_T_411; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_413 = _decoder_T_91 ? 3'h4 : _decoder_T_412; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_414 = _decoder_T_89 ? 3'h2 : _decoder_T_413; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_415 = _decoder_T_87 ? 3'h4 : _decoder_T_414; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_416 = _decoder_T_85 ? 3'h3 : _decoder_T_415; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_417 = _decoder_T_83 ? 3'h4 : _decoder_T_416; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_418 = _decoder_T_75 ? 3'h3 : _decoder_T_417; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_419 = _decoder_T_71 ? 3'h3 : _decoder_T_418; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_420 = _decoder_T_77 ? 3'h4 : _decoder_T_419; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_421 = _decoder_T_75 ? 3'h4 : _decoder_T_420; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_422 = _decoder_T_73 ? 3'h4 : _decoder_T_421; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_423 = _decoder_T_71 ? 3'h4 : _decoder_T_422; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_424 = _decoder_T_69 ? 3'h4 : _decoder_T_423; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_425 = _decoder_T_67 ? 3'h4 : _decoder_T_424; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_426 = _decoder_T_65 ? 3'h2 : _decoder_T_425; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_427 = _decoder_T_63 ? 3'h2 : _decoder_T_426; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_428 = _decoder_T_61 ? 3'h2 : _decoder_T_427; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_429 = _decoder_T_59 ? 3'h2 : _decoder_T_428; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_430 = _decoder_T_57 ? 3'h2 : _decoder_T_429; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_431 = _decoder_T_55 ? 3'h2 : _decoder_T_430; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_432 = _decoder_T_53 ? 3'h1 : _decoder_T_431; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_433 = _decoder_T_51 ? 3'h2 : _decoder_T_432; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_434 = _decoder_T_49 ? 3'h1 : _decoder_T_433; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_435 = _decoder_T_47 ? 3'h2 : _decoder_T_434; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_436 = _decoder_T_45 ? 3'h2 : _decoder_T_435; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_437 = _decoder_T_43 ? 3'h1 : _decoder_T_436; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_438 = _decoder_T_41 ? 3'h1 : _decoder_T_437; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_439 = _decoder_T_39 ? 3'h2 : _decoder_T_438; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_440 = _decoder_T_37 ? 3'h4 : _decoder_T_439; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_441 = _decoder_T_35 ? 3'h4 : _decoder_T_440; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_442 = _decoder_T_33 ? 3'h2 : _decoder_T_441; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_443 = _decoder_T_31 ? 3'h2 : _decoder_T_442; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_444 = _decoder_T_29 ? 3'h4 : _decoder_T_443; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_445 = _decoder_T_27 ? 3'h4 : _decoder_T_444; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_446 = _decoder_T_25 ? 3'h4 : _decoder_T_445; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_447 = _decoder_T_23 ? 3'h4 : _decoder_T_446; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_448 = _decoder_T_21 ? 3'h2 : _decoder_T_447; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_449 = _decoder_T_19 ? 3'h1 : _decoder_T_448; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_450 = _decoder_T_17 ? 3'h2 : _decoder_T_449; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_451 = _decoder_T_15 ? 3'h1 : _decoder_T_450; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_452 = _decoder_T_13 ? 3'h2 : _decoder_T_451; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_453 = _decoder_T_11 ? 3'h2 : _decoder_T_452; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_454 = _decoder_T_9 ? 3'h2 : _decoder_T_453; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_455 = _decoder_T_7 ? 3'h1 : _decoder_T_454; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_456 = _decoder_T_5 ? 3'h2 : _decoder_T_455; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_457 = _decoder_T_3 ? 3'h1 : _decoder_T_456; // @[Lookup.scala 33:37]
  wire [2:0] decoder_5 = _decoder_T_1 ? 3'h2 : _decoder_T_457; // @[Lookup.scala 33:37]
  wire  _decoder_T_475 = _decoder_T_75 ? 1'h0 : _decoder_T_83 | (_decoder_T_85 | (_decoder_T_87 | (_decoder_T_89 | (
    _decoder_T_91 | (_decoder_T_93 | _decoder_T_95))))); // @[Lookup.scala 33:37]
  wire  _decoder_T_476 = _decoder_T_71 ? 1'h0 : _decoder_T_475; // @[Lookup.scala 33:37]
  wire  _decoder_T_477 = _decoder_T_77 ? 1'h0 : _decoder_T_476; // @[Lookup.scala 33:37]
  wire  _decoder_T_478 = _decoder_T_75 ? 1'h0 : _decoder_T_477; // @[Lookup.scala 33:37]
  wire  _decoder_T_479 = _decoder_T_73 ? 1'h0 : _decoder_T_478; // @[Lookup.scala 33:37]
  wire  _decoder_T_480 = _decoder_T_71 ? 1'h0 : _decoder_T_479; // @[Lookup.scala 33:37]
  wire  _decoder_T_481 = _decoder_T_69 ? 1'h0 : _decoder_T_480; // @[Lookup.scala 33:37]
  wire  _decoder_T_482 = _decoder_T_67 ? 1'h0 : _decoder_T_481; // @[Lookup.scala 33:37]
  wire  _decoder_T_483 = _decoder_T_65 ? 1'h0 : _decoder_T_482; // @[Lookup.scala 33:37]
  wire  _decoder_T_484 = _decoder_T_63 ? 1'h0 : _decoder_T_483; // @[Lookup.scala 33:37]
  wire  _decoder_T_485 = _decoder_T_61 ? 1'h0 : _decoder_T_484; // @[Lookup.scala 33:37]
  wire  _decoder_T_486 = _decoder_T_59 ? 1'h0 : _decoder_T_485; // @[Lookup.scala 33:37]
  wire  _decoder_T_487 = _decoder_T_57 ? 1'h0 : _decoder_T_486; // @[Lookup.scala 33:37]
  wire  _decoder_T_488 = _decoder_T_55 ? 1'h0 : _decoder_T_487; // @[Lookup.scala 33:37]
  wire  _decoder_T_489 = _decoder_T_53 ? 1'h0 : _decoder_T_488; // @[Lookup.scala 33:37]
  wire  _decoder_T_490 = _decoder_T_51 ? 1'h0 : _decoder_T_489; // @[Lookup.scala 33:37]
  wire  _decoder_T_491 = _decoder_T_49 ? 1'h0 : _decoder_T_490; // @[Lookup.scala 33:37]
  wire  _decoder_T_492 = _decoder_T_47 ? 1'h0 : _decoder_T_491; // @[Lookup.scala 33:37]
  wire  _decoder_T_493 = _decoder_T_45 ? 1'h0 : _decoder_T_492; // @[Lookup.scala 33:37]
  wire  _decoder_T_494 = _decoder_T_43 ? 1'h0 : _decoder_T_493; // @[Lookup.scala 33:37]
  wire  _decoder_T_495 = _decoder_T_41 ? 1'h0 : _decoder_T_494; // @[Lookup.scala 33:37]
  wire  _decoder_T_496 = _decoder_T_39 ? 1'h0 : _decoder_T_495; // @[Lookup.scala 33:37]
  wire  _decoder_T_497 = _decoder_T_37 ? 1'h0 : _decoder_T_496; // @[Lookup.scala 33:37]
  wire  _decoder_T_498 = _decoder_T_35 ? 1'h0 : _decoder_T_497; // @[Lookup.scala 33:37]
  wire  _decoder_T_499 = _decoder_T_33 ? 1'h0 : _decoder_T_498; // @[Lookup.scala 33:37]
  wire  _decoder_T_500 = _decoder_T_31 ? 1'h0 : _decoder_T_499; // @[Lookup.scala 33:37]
  wire  _decoder_T_501 = _decoder_T_29 ? 1'h0 : _decoder_T_500; // @[Lookup.scala 33:37]
  wire  _decoder_T_502 = _decoder_T_27 ? 1'h0 : _decoder_T_501; // @[Lookup.scala 33:37]
  wire  _decoder_T_503 = _decoder_T_25 ? 1'h0 : _decoder_T_502; // @[Lookup.scala 33:37]
  wire  _decoder_T_504 = _decoder_T_23 ? 1'h0 : _decoder_T_503; // @[Lookup.scala 33:37]
  wire  _decoder_T_505 = _decoder_T_21 ? 1'h0 : _decoder_T_504; // @[Lookup.scala 33:37]
  wire  _decoder_T_506 = _decoder_T_19 ? 1'h0 : _decoder_T_505; // @[Lookup.scala 33:37]
  wire  _decoder_T_507 = _decoder_T_17 ? 1'h0 : _decoder_T_506; // @[Lookup.scala 33:37]
  wire  _decoder_T_508 = _decoder_T_15 ? 1'h0 : _decoder_T_507; // @[Lookup.scala 33:37]
  wire  _decoder_T_509 = _decoder_T_13 ? 1'h0 : _decoder_T_508; // @[Lookup.scala 33:37]
  wire  _decoder_T_510 = _decoder_T_11 ? 1'h0 : _decoder_T_509; // @[Lookup.scala 33:37]
  wire  _decoder_T_511 = _decoder_T_9 ? 1'h0 : _decoder_T_510; // @[Lookup.scala 33:37]
  wire  _decoder_T_512 = _decoder_T_7 ? 1'h0 : _decoder_T_511; // @[Lookup.scala 33:37]
  wire  _decoder_T_513 = _decoder_T_5 ? 1'h0 : _decoder_T_512; // @[Lookup.scala 33:37]
  wire [4:0] rs = io_fb_inst_bank_bits_data_0_inst[25:21]; // @[Decode.scala 34:27]
  wire [4:0] rt = io_fb_inst_bank_bits_data_0_inst[20:16]; // @[Decode.scala 35:27]
  wire [4:0] rd = io_fb_inst_bank_bits_data_0_inst[15:11]; // @[Decode.scala 36:27]
  wire [15:0] rename_info_0_imm_data_lo = io_fb_inst_bank_bits_data_0_inst[15:0]; // @[Decode.scala 37:27]
  wire [25:0] rename_info_0_imm_data_lo_1 = io_fb_inst_bank_bits_data_0_inst[25:0]; // @[Decode.scala 38:27]
  wire [4:0] rename_info_0_imm_data_lo_2 = io_fb_inst_bank_bits_data_0_inst[10:6]; // @[Decode.scala 39:27]
  wire  rename_info_0_need_imm = decoder_2 != 3'h4; // @[Decode.scala 46:25]
  wire [4:0] _rename_info_0_op1_addr_T_6 = 3'h0 == decoder_3 ? rs : 5'h0; // @[Mux.scala 80:57]
  wire [4:0] _rename_info_0_op1_addr_T_8 = 3'h1 == decoder_3 ? rt : _rename_info_0_op1_addr_T_6; // @[Mux.scala 80:57]
  wire [4:0] _rename_info_0_op1_addr_T_10 = 3'h2 == decoder_3 ? rd : _rename_info_0_op1_addr_T_8; // @[Mux.scala 80:57]
  wire [4:0] rename_info_0_op1_addr = 3'h3 == decoder_3 ? 5'h1f : _rename_info_0_op1_addr_T_10; // @[Mux.scala 80:57]
  wire [4:0] _rename_info_0_op2_addr_T_6 = 3'h0 == decoder_4 ? rs : 5'h0; // @[Mux.scala 80:57]
  wire [4:0] _rename_info_0_op2_addr_T_8 = 3'h1 == decoder_4 ? rt : _rename_info_0_op2_addr_T_6; // @[Mux.scala 80:57]
  wire [4:0] _rename_info_0_op2_addr_T_10 = 3'h2 == decoder_4 ? rd : _rename_info_0_op2_addr_T_8; // @[Mux.scala 80:57]
  wire [4:0] rename_info_0_op2_addr = 3'h3 == decoder_4 ? 5'h1f : _rename_info_0_op2_addr_T_10; // @[Mux.scala 80:57]
  wire [4:0] _rename_info_0_des_addr_T_6 = 3'h0 == decoder_5 ? rs : 5'h0; // @[Mux.scala 80:57]
  wire [4:0] _rename_info_0_des_addr_T_8 = 3'h1 == decoder_5 ? rt : _rename_info_0_des_addr_T_6; // @[Mux.scala 80:57]
  wire [4:0] _rename_info_0_des_addr_T_10 = 3'h2 == decoder_5 ? rd : _rename_info_0_des_addr_T_8; // @[Mux.scala 80:57]
  wire [4:0] rename_info_0_des_addr = 3'h3 == decoder_5 ? 5'h1f : _rename_info_0_des_addr_T_10; // @[Mux.scala 80:57]
  wire [15:0] rename_info_0_imm_data_hi = rename_info_0_imm_data_lo[15] ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _rename_info_0_imm_data_T_4 = {rename_info_0_imm_data_hi,rename_info_0_imm_data_lo}; // @[Cat.scala 30:58]
  wire [31:0] _rename_info_0_imm_data_T_6 = {16'h0,rename_info_0_imm_data_lo}; // @[Cat.scala 30:58]
  wire [31:0] _rename_info_0_imm_data_T_8 = {27'h0,rename_info_0_imm_data_lo_2}; // @[Cat.scala 30:58]
  wire [35:0] _rename_info_0_imm_data_T_10 = {10'h0,rename_info_0_imm_data_lo_1}; // @[Cat.scala 30:58]
  wire [31:0] _rename_info_0_imm_data_T_12 = 3'h1 == decoder_2 ? _rename_info_0_imm_data_T_4 : 32'h0; // @[Mux.scala 80:57]
  wire [31:0] _rename_info_0_imm_data_T_14 = 3'h0 == decoder_2 ? _rename_info_0_imm_data_T_6 :
    _rename_info_0_imm_data_T_12; // @[Mux.scala 80:57]
  wire [31:0] _rename_info_0_imm_data_T_16 = 3'h2 == decoder_2 ? _rename_info_0_imm_data_T_8 :
    _rename_info_0_imm_data_T_14; // @[Mux.scala 80:57]
  wire [35:0] _rename_info_0_imm_data_T_18 = 3'h3 == decoder_2 ? _rename_info_0_imm_data_T_10 : {{4'd0},
    _rename_info_0_imm_data_T_16}; // @[Mux.scala 80:57]
  wire [31:0] _decoder_T_572 = io_fb_inst_bank_bits_data_1_inst & 32'hfc0007ff; // @[Lookup.scala 31:38]
  wire  _decoder_T_573 = 32'h20 == _decoder_T_572; // @[Lookup.scala 31:38]
  wire [31:0] _decoder_T_574 = io_fb_inst_bank_bits_data_1_inst & 32'hfc000000; // @[Lookup.scala 31:38]
  wire  _decoder_T_575 = 32'h20000000 == _decoder_T_574; // @[Lookup.scala 31:38]
  wire  _decoder_T_577 = 32'h21 == _decoder_T_572; // @[Lookup.scala 31:38]
  wire  _decoder_T_579 = 32'h24000000 == _decoder_T_574; // @[Lookup.scala 31:38]
  wire  _decoder_T_581 = 32'h22 == _decoder_T_572; // @[Lookup.scala 31:38]
  wire  _decoder_T_583 = 32'h23 == _decoder_T_572; // @[Lookup.scala 31:38]
  wire  _decoder_T_585 = 32'h2a == _decoder_T_572; // @[Lookup.scala 31:38]
  wire  _decoder_T_587 = 32'h28000000 == _decoder_T_574; // @[Lookup.scala 31:38]
  wire  _decoder_T_589 = 32'h2b == _decoder_T_572; // @[Lookup.scala 31:38]
  wire  _decoder_T_591 = 32'h2c000000 == _decoder_T_574; // @[Lookup.scala 31:38]
  wire  _decoder_T_593 = 32'h70000002 == _decoder_T_572; // @[Lookup.scala 31:38]
  wire [31:0] _decoder_T_594 = io_fb_inst_bank_bits_data_1_inst & 32'hfc00ffff; // @[Lookup.scala 31:38]
  wire  _decoder_T_595 = 32'h1a == _decoder_T_594; // @[Lookup.scala 31:38]
  wire  _decoder_T_597 = 32'h1b == _decoder_T_594; // @[Lookup.scala 31:38]
  wire  _decoder_T_599 = 32'h18 == _decoder_T_594; // @[Lookup.scala 31:38]
  wire  _decoder_T_601 = 32'h19 == _decoder_T_594; // @[Lookup.scala 31:38]
  wire [31:0] _decoder_T_602 = io_fb_inst_bank_bits_data_1_inst & 32'hffff07ff; // @[Lookup.scala 31:38]
  wire  _decoder_T_603 = 32'h10 == _decoder_T_602; // @[Lookup.scala 31:38]
  wire  _decoder_T_605 = 32'h12 == _decoder_T_602; // @[Lookup.scala 31:38]
  wire [31:0] _decoder_T_606 = io_fb_inst_bank_bits_data_1_inst & 32'hfc1fffff; // @[Lookup.scala 31:38]
  wire  _decoder_T_607 = 32'h11 == _decoder_T_606; // @[Lookup.scala 31:38]
  wire  _decoder_T_609 = 32'h13 == _decoder_T_606; // @[Lookup.scala 31:38]
  wire  _decoder_T_611 = 32'h24 == _decoder_T_572; // @[Lookup.scala 31:38]
  wire  _decoder_T_613 = 32'h30000000 == _decoder_T_574; // @[Lookup.scala 31:38]
  wire [31:0] _decoder_T_614 = io_fb_inst_bank_bits_data_1_inst & 32'hffe00000; // @[Lookup.scala 31:38]
  wire  _decoder_T_615 = 32'h3c000000 == _decoder_T_614; // @[Lookup.scala 31:38]
  wire  _decoder_T_617 = 32'h27 == _decoder_T_572; // @[Lookup.scala 31:38]
  wire  _decoder_T_619 = 32'h25 == _decoder_T_572; // @[Lookup.scala 31:38]
  wire  _decoder_T_621 = 32'h34000000 == _decoder_T_574; // @[Lookup.scala 31:38]
  wire  _decoder_T_623 = 32'h26 == _decoder_T_572; // @[Lookup.scala 31:38]
  wire  _decoder_T_625 = 32'h38000000 == _decoder_T_574; // @[Lookup.scala 31:38]
  wire  _decoder_T_627 = 32'h4 == _decoder_T_572; // @[Lookup.scala 31:38]
  wire [31:0] _decoder_T_628 = io_fb_inst_bank_bits_data_1_inst & 32'hffe0003f; // @[Lookup.scala 31:38]
  wire  _decoder_T_629 = 32'h0 == _decoder_T_628; // @[Lookup.scala 31:38]
  wire  _decoder_T_631 = 32'h7 == _decoder_T_572; // @[Lookup.scala 31:38]
  wire  _decoder_T_633 = 32'h3 == _decoder_T_628; // @[Lookup.scala 31:38]
  wire  _decoder_T_635 = 32'h6 == _decoder_T_572; // @[Lookup.scala 31:38]
  wire  _decoder_T_637 = 32'h2 == _decoder_T_628; // @[Lookup.scala 31:38]
  wire  _decoder_T_639 = 32'h10000000 == _decoder_T_574; // @[Lookup.scala 31:38]
  wire  _decoder_T_641 = 32'h14000000 == _decoder_T_574; // @[Lookup.scala 31:38]
  wire [31:0] _decoder_T_642 = io_fb_inst_bank_bits_data_1_inst & 32'hfc1f0000; // @[Lookup.scala 31:38]
  wire  _decoder_T_643 = 32'h4010000 == _decoder_T_642; // @[Lookup.scala 31:38]
  wire  _decoder_T_645 = 32'h1c000000 == _decoder_T_642; // @[Lookup.scala 31:38]
  wire  _decoder_T_647 = 32'h18000000 == _decoder_T_642; // @[Lookup.scala 31:38]
  wire  _decoder_T_649 = 32'h4000000 == _decoder_T_642; // @[Lookup.scala 31:38]
  wire  _decoder_T_655 = 32'h8000000 == _decoder_T_574; // @[Lookup.scala 31:38]
  wire  _decoder_T_657 = 32'hc000000 == _decoder_T_574; // @[Lookup.scala 31:38]
  wire  _decoder_T_659 = 32'h8 == _decoder_T_606; // @[Lookup.scala 31:38]
  wire [31:0] _decoder_T_660 = io_fb_inst_bank_bits_data_1_inst & 32'hfc1f07ff; // @[Lookup.scala 31:38]
  wire  _decoder_T_661 = 32'h9 == _decoder_T_660; // @[Lookup.scala 31:38]
  wire  _decoder_T_663 = 32'hc == io_fb_inst_bank_bits_data_1_inst; // @[Lookup.scala 31:38]
  wire [31:0] _decoder_T_664 = io_fb_inst_bank_bits_data_1_inst & 32'hfc00003f; // @[Lookup.scala 31:38]
  wire  _decoder_T_665 = 32'hd == _decoder_T_664; // @[Lookup.scala 31:38]
  wire  _decoder_T_667 = 32'h42000018 == io_fb_inst_bank_bits_data_1_inst; // @[Lookup.scala 31:38]
  wire [31:0] _decoder_T_668 = io_fb_inst_bank_bits_data_1_inst & 32'hffe007ff; // @[Lookup.scala 31:38]
  wire  _decoder_T_669 = 32'h40000000 == _decoder_T_668; // @[Lookup.scala 31:38]
  wire  _decoder_T_671 = 32'h40800000 == _decoder_T_668; // @[Lookup.scala 31:38]
  wire  _decoder_T_673 = 32'h80000000 == _decoder_T_574; // @[Lookup.scala 31:38]
  wire  _decoder_T_675 = 32'h84000000 == _decoder_T_574; // @[Lookup.scala 31:38]
  wire  _decoder_T_677 = 32'h8c000000 == _decoder_T_574; // @[Lookup.scala 31:38]
  wire  _decoder_T_679 = 32'h90000000 == _decoder_T_574; // @[Lookup.scala 31:38]
  wire  _decoder_T_681 = 32'h94000000 == _decoder_T_574; // @[Lookup.scala 31:38]
  wire  _decoder_T_683 = 32'ha0000000 == _decoder_T_574; // @[Lookup.scala 31:38]
  wire  _decoder_T_685 = 32'ha4000000 == _decoder_T_574; // @[Lookup.scala 31:38]
  wire  _decoder_T_687 = 32'hac000000 == _decoder_T_574; // @[Lookup.scala 31:38]
  wire [5:0] _decoder_T_688 = _decoder_T_687 ? 6'h24 : 6'h0; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_689 = _decoder_T_685 ? 6'h25 : _decoder_T_688; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_690 = _decoder_T_683 ? 6'h26 : _decoder_T_689; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_691 = _decoder_T_681 ? 6'h29 : _decoder_T_690; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_692 = _decoder_T_679 ? 6'h2b : _decoder_T_691; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_693 = _decoder_T_677 ? 6'h27 : _decoder_T_692; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_694 = _decoder_T_675 ? 6'h28 : _decoder_T_693; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_695 = _decoder_T_673 ? 6'h2a : _decoder_T_694; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_696 = _decoder_T_671 ? 6'h2c : _decoder_T_695; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_697 = _decoder_T_669 ? 6'h2d : _decoder_T_696; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_698 = _decoder_T_667 ? 6'h2f : _decoder_T_697; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_699 = _decoder_T_665 ? 6'h30 : _decoder_T_698; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_700 = _decoder_T_663 ? 6'h2e : _decoder_T_699; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_701 = _decoder_T_661 ? 6'h1b : _decoder_T_700; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_702 = _decoder_T_659 ? 6'h1a : _decoder_T_701; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_703 = _decoder_T_657 ? 6'h19 : _decoder_T_702; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_704 = _decoder_T_655 ? 6'h18 : _decoder_T_703; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_705 = _decoder_T_647 ? 6'h23 : _decoder_T_704; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_706 = _decoder_T_643 ? 6'h22 : _decoder_T_705; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_707 = _decoder_T_649 ? 6'h20 : _decoder_T_706; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_708 = _decoder_T_647 ? 6'h1e : _decoder_T_707; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_709 = _decoder_T_645 ? 6'h1f : _decoder_T_708; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_710 = _decoder_T_643 ? 6'h21 : _decoder_T_709; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_711 = _decoder_T_641 ? 6'h1d : _decoder_T_710; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_712 = _decoder_T_639 ? 6'h1c : _decoder_T_711; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_713 = _decoder_T_637 ? 6'h6 : _decoder_T_712; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_714 = _decoder_T_635 ? 6'h6 : _decoder_T_713; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_715 = _decoder_T_633 ? 6'h7 : _decoder_T_714; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_716 = _decoder_T_631 ? 6'h7 : _decoder_T_715; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_717 = _decoder_T_629 ? 6'h5 : _decoder_T_716; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_718 = _decoder_T_627 ? 6'h5 : _decoder_T_717; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_719 = _decoder_T_625 ? 6'ha : _decoder_T_718; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_720 = _decoder_T_623 ? 6'ha : _decoder_T_719; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_721 = _decoder_T_621 ? 6'hb : _decoder_T_720; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_722 = _decoder_T_619 ? 6'hb : _decoder_T_721; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_723 = _decoder_T_617 ? 6'he : _decoder_T_722; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_724 = _decoder_T_615 ? 6'hd : _decoder_T_723; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_725 = _decoder_T_613 ? 6'hc : _decoder_T_724; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_726 = _decoder_T_611 ? 6'hc : _decoder_T_725; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_727 = _decoder_T_609 ? 6'h17 : _decoder_T_726; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_728 = _decoder_T_607 ? 6'h16 : _decoder_T_727; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_729 = _decoder_T_605 ? 6'h15 : _decoder_T_728; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_730 = _decoder_T_603 ? 6'h14 : _decoder_T_729; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_731 = _decoder_T_601 ? 6'h11 : _decoder_T_730; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_732 = _decoder_T_599 ? 6'h10 : _decoder_T_731; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_733 = _decoder_T_597 ? 6'h13 : _decoder_T_732; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_734 = _decoder_T_595 ? 6'h12 : _decoder_T_733; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_735 = _decoder_T_593 ? 6'hf : _decoder_T_734; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_736 = _decoder_T_591 ? 6'h9 : _decoder_T_735; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_737 = _decoder_T_589 ? 6'h9 : _decoder_T_736; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_738 = _decoder_T_587 ? 6'h8 : _decoder_T_737; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_739 = _decoder_T_585 ? 6'h8 : _decoder_T_738; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_740 = _decoder_T_583 ? 6'h4 : _decoder_T_739; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_741 = _decoder_T_581 ? 6'h3 : _decoder_T_740; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_742 = _decoder_T_579 ? 6'h2 : _decoder_T_741; // @[Lookup.scala 33:37]
  wire [5:0] _decoder_T_743 = _decoder_T_577 ? 6'h2 : _decoder_T_742; // @[Lookup.scala 33:37]
  wire [1:0] _decoder_T_745 = _decoder_T_687 ? 2'h3 : 2'h0; // @[Lookup.scala 33:37]
  wire [1:0] _decoder_T_746 = _decoder_T_685 ? 2'h3 : _decoder_T_745; // @[Lookup.scala 33:37]
  wire [1:0] _decoder_T_747 = _decoder_T_683 ? 2'h3 : _decoder_T_746; // @[Lookup.scala 33:37]
  wire [1:0] _decoder_T_748 = _decoder_T_681 ? 2'h3 : _decoder_T_747; // @[Lookup.scala 33:37]
  wire [1:0] _decoder_T_749 = _decoder_T_679 ? 2'h3 : _decoder_T_748; // @[Lookup.scala 33:37]
  wire [1:0] _decoder_T_750 = _decoder_T_677 ? 2'h3 : _decoder_T_749; // @[Lookup.scala 33:37]
  wire [1:0] _decoder_T_751 = _decoder_T_675 ? 2'h3 : _decoder_T_750; // @[Lookup.scala 33:37]
  wire [1:0] _decoder_T_752 = _decoder_T_673 ? 2'h3 : _decoder_T_751; // @[Lookup.scala 33:37]
  wire [1:0] _decoder_T_753 = _decoder_T_671 ? 2'h2 : _decoder_T_752; // @[Lookup.scala 33:37]
  wire [1:0] _decoder_T_754 = _decoder_T_669 ? 2'h2 : _decoder_T_753; // @[Lookup.scala 33:37]
  wire [1:0] _decoder_T_755 = _decoder_T_667 ? 2'h0 : _decoder_T_754; // @[Lookup.scala 33:37]
  wire [1:0] _decoder_T_756 = _decoder_T_665 ? 2'h0 : _decoder_T_755; // @[Lookup.scala 33:37]
  wire [1:0] _decoder_T_757 = _decoder_T_663 ? 2'h0 : _decoder_T_756; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_758 = _decoder_T_661 ? 3'h5 : {{1'd0}, _decoder_T_757}; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_759 = _decoder_T_659 ? 3'h5 : _decoder_T_758; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_760 = _decoder_T_657 ? 3'h5 : _decoder_T_759; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_761 = _decoder_T_655 ? 3'h5 : _decoder_T_760; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_762 = _decoder_T_647 ? 3'h5 : _decoder_T_761; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_763 = _decoder_T_643 ? 3'h5 : _decoder_T_762; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_764 = _decoder_T_649 ? 3'h5 : _decoder_T_763; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_765 = _decoder_T_647 ? 3'h5 : _decoder_T_764; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_766 = _decoder_T_645 ? 3'h5 : _decoder_T_765; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_767 = _decoder_T_643 ? 3'h5 : _decoder_T_766; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_768 = _decoder_T_641 ? 3'h5 : _decoder_T_767; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_769 = _decoder_T_639 ? 3'h5 : _decoder_T_768; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_770 = _decoder_T_637 ? 3'h1 : _decoder_T_769; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_771 = _decoder_T_635 ? 3'h1 : _decoder_T_770; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_772 = _decoder_T_633 ? 3'h1 : _decoder_T_771; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_773 = _decoder_T_631 ? 3'h1 : _decoder_T_772; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_774 = _decoder_T_629 ? 3'h1 : _decoder_T_773; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_775 = _decoder_T_627 ? 3'h1 : _decoder_T_774; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_776 = _decoder_T_625 ? 3'h1 : _decoder_T_775; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_777 = _decoder_T_623 ? 3'h1 : _decoder_T_776; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_778 = _decoder_T_621 ? 3'h1 : _decoder_T_777; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_779 = _decoder_T_619 ? 3'h1 : _decoder_T_778; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_780 = _decoder_T_617 ? 3'h1 : _decoder_T_779; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_781 = _decoder_T_615 ? 3'h1 : _decoder_T_780; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_782 = _decoder_T_613 ? 3'h1 : _decoder_T_781; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_783 = _decoder_T_611 ? 3'h1 : _decoder_T_782; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_784 = _decoder_T_609 ? 3'h4 : _decoder_T_783; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_785 = _decoder_T_607 ? 3'h4 : _decoder_T_784; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_786 = _decoder_T_605 ? 3'h4 : _decoder_T_785; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_787 = _decoder_T_603 ? 3'h4 : _decoder_T_786; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_788 = _decoder_T_601 ? 3'h4 : _decoder_T_787; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_789 = _decoder_T_599 ? 3'h4 : _decoder_T_788; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_790 = _decoder_T_597 ? 3'h4 : _decoder_T_789; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_791 = _decoder_T_595 ? 3'h4 : _decoder_T_790; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_792 = _decoder_T_593 ? 3'h4 : _decoder_T_791; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_793 = _decoder_T_591 ? 3'h1 : _decoder_T_792; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_794 = _decoder_T_589 ? 3'h1 : _decoder_T_793; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_795 = _decoder_T_587 ? 3'h1 : _decoder_T_794; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_796 = _decoder_T_585 ? 3'h1 : _decoder_T_795; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_797 = _decoder_T_583 ? 3'h1 : _decoder_T_796; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_798 = _decoder_T_581 ? 3'h1 : _decoder_T_797; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_799 = _decoder_T_579 ? 3'h1 : _decoder_T_798; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_800 = _decoder_T_577 ? 3'h1 : _decoder_T_799; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_802 = _decoder_T_687 ? 3'h1 : 3'h4; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_803 = _decoder_T_685 ? 3'h1 : _decoder_T_802; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_804 = _decoder_T_683 ? 3'h1 : _decoder_T_803; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_805 = _decoder_T_681 ? 3'h1 : _decoder_T_804; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_806 = _decoder_T_679 ? 3'h1 : _decoder_T_805; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_807 = _decoder_T_677 ? 3'h1 : _decoder_T_806; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_808 = _decoder_T_675 ? 3'h1 : _decoder_T_807; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_809 = _decoder_T_673 ? 3'h1 : _decoder_T_808; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_810 = _decoder_T_671 ? 3'h0 : _decoder_T_809; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_811 = _decoder_T_669 ? 3'h0 : _decoder_T_810; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_812 = _decoder_T_667 ? 3'h4 : _decoder_T_811; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_813 = _decoder_T_665 ? 3'h4 : _decoder_T_812; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_814 = _decoder_T_663 ? 3'h4 : _decoder_T_813; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_815 = _decoder_T_661 ? 3'h4 : _decoder_T_814; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_816 = _decoder_T_659 ? 3'h4 : _decoder_T_815; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_817 = _decoder_T_657 ? 3'h3 : _decoder_T_816; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_818 = _decoder_T_655 ? 3'h3 : _decoder_T_817; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_819 = _decoder_T_647 ? 3'h1 : _decoder_T_818; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_820 = _decoder_T_643 ? 3'h1 : _decoder_T_819; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_821 = _decoder_T_649 ? 3'h1 : _decoder_T_820; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_822 = _decoder_T_647 ? 3'h1 : _decoder_T_821; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_823 = _decoder_T_645 ? 3'h1 : _decoder_T_822; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_824 = _decoder_T_643 ? 3'h1 : _decoder_T_823; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_825 = _decoder_T_641 ? 3'h1 : _decoder_T_824; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_826 = _decoder_T_639 ? 3'h1 : _decoder_T_825; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_827 = _decoder_T_637 ? 3'h2 : _decoder_T_826; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_828 = _decoder_T_635 ? 3'h4 : _decoder_T_827; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_829 = _decoder_T_633 ? 3'h2 : _decoder_T_828; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_830 = _decoder_T_631 ? 3'h4 : _decoder_T_829; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_831 = _decoder_T_629 ? 3'h2 : _decoder_T_830; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_832 = _decoder_T_627 ? 3'h4 : _decoder_T_831; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_833 = _decoder_T_625 ? 3'h0 : _decoder_T_832; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_834 = _decoder_T_623 ? 3'h4 : _decoder_T_833; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_835 = _decoder_T_621 ? 3'h0 : _decoder_T_834; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_836 = _decoder_T_619 ? 3'h4 : _decoder_T_835; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_837 = _decoder_T_617 ? 3'h4 : _decoder_T_836; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_838 = _decoder_T_615 ? 3'h0 : _decoder_T_837; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_839 = _decoder_T_613 ? 3'h0 : _decoder_T_838; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_840 = _decoder_T_611 ? 3'h4 : _decoder_T_839; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_841 = _decoder_T_609 ? 3'h4 : _decoder_T_840; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_842 = _decoder_T_607 ? 3'h4 : _decoder_T_841; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_843 = _decoder_T_605 ? 3'h4 : _decoder_T_842; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_844 = _decoder_T_603 ? 3'h4 : _decoder_T_843; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_845 = _decoder_T_601 ? 3'h4 : _decoder_T_844; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_846 = _decoder_T_599 ? 3'h4 : _decoder_T_845; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_847 = _decoder_T_597 ? 3'h4 : _decoder_T_846; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_848 = _decoder_T_595 ? 3'h4 : _decoder_T_847; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_849 = _decoder_T_593 ? 3'h4 : _decoder_T_848; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_850 = _decoder_T_591 ? 3'h1 : _decoder_T_849; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_851 = _decoder_T_589 ? 3'h4 : _decoder_T_850; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_852 = _decoder_T_587 ? 3'h1 : _decoder_T_851; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_853 = _decoder_T_585 ? 3'h4 : _decoder_T_852; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_854 = _decoder_T_583 ? 3'h4 : _decoder_T_853; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_855 = _decoder_T_581 ? 3'h4 : _decoder_T_854; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_856 = _decoder_T_579 ? 3'h1 : _decoder_T_855; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_857 = _decoder_T_577 ? 3'h4 : _decoder_T_856; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_858 = _decoder_T_575 ? 3'h1 : _decoder_T_857; // @[Lookup.scala 33:37]
  wire [2:0] decoder_2_1 = _decoder_T_573 ? 3'h4 : _decoder_T_858; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_859 = _decoder_T_687 ? 3'h0 : 3'h4; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_860 = _decoder_T_685 ? 3'h0 : _decoder_T_859; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_861 = _decoder_T_683 ? 3'h0 : _decoder_T_860; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_862 = _decoder_T_681 ? 3'h0 : _decoder_T_861; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_863 = _decoder_T_679 ? 3'h0 : _decoder_T_862; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_864 = _decoder_T_677 ? 3'h0 : _decoder_T_863; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_865 = _decoder_T_675 ? 3'h0 : _decoder_T_864; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_866 = _decoder_T_673 ? 3'h0 : _decoder_T_865; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_867 = _decoder_T_671 ? 3'h1 : _decoder_T_866; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_868 = _decoder_T_669 ? 3'h2 : _decoder_T_867; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_869 = _decoder_T_667 ? 3'h4 : _decoder_T_868; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_870 = _decoder_T_665 ? 3'h4 : _decoder_T_869; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_871 = _decoder_T_663 ? 3'h4 : _decoder_T_870; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_872 = _decoder_T_661 ? 3'h0 : _decoder_T_871; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_873 = _decoder_T_659 ? 3'h0 : _decoder_T_872; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_874 = _decoder_T_657 ? 3'h4 : _decoder_T_873; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_875 = _decoder_T_655 ? 3'h4 : _decoder_T_874; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_876 = _decoder_T_647 ? 3'h0 : _decoder_T_875; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_877 = _decoder_T_643 ? 3'h0 : _decoder_T_876; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_878 = _decoder_T_649 ? 3'h0 : _decoder_T_877; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_879 = _decoder_T_647 ? 3'h0 : _decoder_T_878; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_880 = _decoder_T_645 ? 3'h0 : _decoder_T_879; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_881 = _decoder_T_643 ? 3'h0 : _decoder_T_880; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_882 = _decoder_T_641 ? 3'h0 : _decoder_T_881; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_883 = _decoder_T_639 ? 3'h0 : _decoder_T_882; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_884 = _decoder_T_637 ? 3'h1 : _decoder_T_883; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_885 = _decoder_T_635 ? 3'h1 : _decoder_T_884; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_886 = _decoder_T_633 ? 3'h1 : _decoder_T_885; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_887 = _decoder_T_631 ? 3'h1 : _decoder_T_886; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_888 = _decoder_T_629 ? 3'h1 : _decoder_T_887; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_889 = _decoder_T_627 ? 3'h1 : _decoder_T_888; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_890 = _decoder_T_625 ? 3'h0 : _decoder_T_889; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_891 = _decoder_T_623 ? 3'h0 : _decoder_T_890; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_892 = _decoder_T_621 ? 3'h0 : _decoder_T_891; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_893 = _decoder_T_619 ? 3'h0 : _decoder_T_892; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_894 = _decoder_T_617 ? 3'h0 : _decoder_T_893; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_895 = _decoder_T_615 ? 3'h4 : _decoder_T_894; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_896 = _decoder_T_613 ? 3'h0 : _decoder_T_895; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_897 = _decoder_T_611 ? 3'h0 : _decoder_T_896; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_898 = _decoder_T_609 ? 3'h0 : _decoder_T_897; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_899 = _decoder_T_607 ? 3'h0 : _decoder_T_898; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_900 = _decoder_T_605 ? 3'h4 : _decoder_T_899; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_901 = _decoder_T_603 ? 3'h4 : _decoder_T_900; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_902 = _decoder_T_601 ? 3'h0 : _decoder_T_901; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_903 = _decoder_T_599 ? 3'h0 : _decoder_T_902; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_904 = _decoder_T_597 ? 3'h0 : _decoder_T_903; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_905 = _decoder_T_595 ? 3'h0 : _decoder_T_904; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_906 = _decoder_T_593 ? 3'h0 : _decoder_T_905; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_907 = _decoder_T_591 ? 3'h0 : _decoder_T_906; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_908 = _decoder_T_589 ? 3'h0 : _decoder_T_907; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_909 = _decoder_T_587 ? 3'h0 : _decoder_T_908; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_910 = _decoder_T_585 ? 3'h0 : _decoder_T_909; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_911 = _decoder_T_583 ? 3'h0 : _decoder_T_910; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_912 = _decoder_T_581 ? 3'h0 : _decoder_T_911; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_913 = _decoder_T_579 ? 3'h0 : _decoder_T_912; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_914 = _decoder_T_577 ? 3'h0 : _decoder_T_913; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_915 = _decoder_T_575 ? 3'h0 : _decoder_T_914; // @[Lookup.scala 33:37]
  wire [2:0] decoder_3_1 = _decoder_T_573 ? 3'h0 : _decoder_T_915; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_919 = _decoder_T_681 ? 3'h4 : _decoder_T_804; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_920 = _decoder_T_679 ? 3'h4 : _decoder_T_919; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_921 = _decoder_T_677 ? 3'h4 : _decoder_T_920; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_922 = _decoder_T_675 ? 3'h4 : _decoder_T_921; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_923 = _decoder_T_673 ? 3'h4 : _decoder_T_922; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_924 = _decoder_T_671 ? 3'h2 : _decoder_T_923; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_925 = _decoder_T_669 ? 3'h4 : _decoder_T_924; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_926 = _decoder_T_667 ? 3'h4 : _decoder_T_925; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_927 = _decoder_T_665 ? 3'h4 : _decoder_T_926; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_928 = _decoder_T_663 ? 3'h4 : _decoder_T_927; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_929 = _decoder_T_661 ? 3'h4 : _decoder_T_928; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_930 = _decoder_T_659 ? 3'h4 : _decoder_T_929; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_931 = _decoder_T_657 ? 3'h4 : _decoder_T_930; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_932 = _decoder_T_655 ? 3'h4 : _decoder_T_931; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_933 = _decoder_T_647 ? 3'h4 : _decoder_T_932; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_934 = _decoder_T_643 ? 3'h4 : _decoder_T_933; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_935 = _decoder_T_649 ? 3'h4 : _decoder_T_934; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_936 = _decoder_T_647 ? 3'h4 : _decoder_T_935; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_937 = _decoder_T_645 ? 3'h4 : _decoder_T_936; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_938 = _decoder_T_643 ? 3'h4 : _decoder_T_937; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_939 = _decoder_T_641 ? 3'h1 : _decoder_T_938; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_940 = _decoder_T_639 ? 3'h1 : _decoder_T_939; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_941 = _decoder_T_637 ? 3'h4 : _decoder_T_940; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_942 = _decoder_T_635 ? 3'h0 : _decoder_T_941; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_943 = _decoder_T_633 ? 3'h4 : _decoder_T_942; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_944 = _decoder_T_631 ? 3'h0 : _decoder_T_943; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_945 = _decoder_T_629 ? 3'h4 : _decoder_T_944; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_946 = _decoder_T_627 ? 3'h0 : _decoder_T_945; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_947 = _decoder_T_625 ? 3'h4 : _decoder_T_946; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_948 = _decoder_T_623 ? 3'h1 : _decoder_T_947; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_949 = _decoder_T_621 ? 3'h4 : _decoder_T_948; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_950 = _decoder_T_619 ? 3'h1 : _decoder_T_949; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_951 = _decoder_T_617 ? 3'h1 : _decoder_T_950; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_952 = _decoder_T_615 ? 3'h4 : _decoder_T_951; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_953 = _decoder_T_613 ? 3'h4 : _decoder_T_952; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_954 = _decoder_T_611 ? 3'h1 : _decoder_T_953; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_955 = _decoder_T_609 ? 3'h4 : _decoder_T_954; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_956 = _decoder_T_607 ? 3'h4 : _decoder_T_955; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_957 = _decoder_T_605 ? 3'h4 : _decoder_T_956; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_958 = _decoder_T_603 ? 3'h4 : _decoder_T_957; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_959 = _decoder_T_601 ? 3'h1 : _decoder_T_958; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_960 = _decoder_T_599 ? 3'h1 : _decoder_T_959; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_961 = _decoder_T_597 ? 3'h1 : _decoder_T_960; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_962 = _decoder_T_595 ? 3'h1 : _decoder_T_961; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_963 = _decoder_T_593 ? 3'h1 : _decoder_T_962; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_964 = _decoder_T_591 ? 3'h4 : _decoder_T_963; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_965 = _decoder_T_589 ? 3'h1 : _decoder_T_964; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_966 = _decoder_T_587 ? 3'h4 : _decoder_T_965; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_967 = _decoder_T_585 ? 3'h1 : _decoder_T_966; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_968 = _decoder_T_583 ? 3'h1 : _decoder_T_967; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_969 = _decoder_T_581 ? 3'h1 : _decoder_T_968; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_970 = _decoder_T_579 ? 3'h4 : _decoder_T_969; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_971 = _decoder_T_577 ? 3'h1 : _decoder_T_970; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_972 = _decoder_T_575 ? 3'h4 : _decoder_T_971; // @[Lookup.scala 33:37]
  wire [2:0] decoder_4_1 = _decoder_T_573 ? 3'h1 : _decoder_T_972; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_976 = _decoder_T_681 ? 3'h1 : 3'h4; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_977 = _decoder_T_679 ? 3'h1 : _decoder_T_976; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_978 = _decoder_T_677 ? 3'h1 : _decoder_T_977; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_979 = _decoder_T_675 ? 3'h1 : _decoder_T_978; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_980 = _decoder_T_673 ? 3'h1 : _decoder_T_979; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_981 = _decoder_T_671 ? 3'h4 : _decoder_T_980; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_982 = _decoder_T_669 ? 3'h1 : _decoder_T_981; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_983 = _decoder_T_667 ? 3'h4 : _decoder_T_982; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_984 = _decoder_T_665 ? 3'h4 : _decoder_T_983; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_985 = _decoder_T_663 ? 3'h4 : _decoder_T_984; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_986 = _decoder_T_661 ? 3'h2 : _decoder_T_985; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_987 = _decoder_T_659 ? 3'h4 : _decoder_T_986; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_988 = _decoder_T_657 ? 3'h3 : _decoder_T_987; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_989 = _decoder_T_655 ? 3'h4 : _decoder_T_988; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_990 = _decoder_T_647 ? 3'h3 : _decoder_T_989; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_991 = _decoder_T_643 ? 3'h3 : _decoder_T_990; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_992 = _decoder_T_649 ? 3'h4 : _decoder_T_991; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_993 = _decoder_T_647 ? 3'h4 : _decoder_T_992; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_994 = _decoder_T_645 ? 3'h4 : _decoder_T_993; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_995 = _decoder_T_643 ? 3'h4 : _decoder_T_994; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_996 = _decoder_T_641 ? 3'h4 : _decoder_T_995; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_997 = _decoder_T_639 ? 3'h4 : _decoder_T_996; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_998 = _decoder_T_637 ? 3'h2 : _decoder_T_997; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_999 = _decoder_T_635 ? 3'h2 : _decoder_T_998; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_1000 = _decoder_T_633 ? 3'h2 : _decoder_T_999; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_1001 = _decoder_T_631 ? 3'h2 : _decoder_T_1000; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_1002 = _decoder_T_629 ? 3'h2 : _decoder_T_1001; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_1003 = _decoder_T_627 ? 3'h2 : _decoder_T_1002; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_1004 = _decoder_T_625 ? 3'h1 : _decoder_T_1003; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_1005 = _decoder_T_623 ? 3'h2 : _decoder_T_1004; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_1006 = _decoder_T_621 ? 3'h1 : _decoder_T_1005; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_1007 = _decoder_T_619 ? 3'h2 : _decoder_T_1006; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_1008 = _decoder_T_617 ? 3'h2 : _decoder_T_1007; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_1009 = _decoder_T_615 ? 3'h1 : _decoder_T_1008; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_1010 = _decoder_T_613 ? 3'h1 : _decoder_T_1009; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_1011 = _decoder_T_611 ? 3'h2 : _decoder_T_1010; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_1012 = _decoder_T_609 ? 3'h4 : _decoder_T_1011; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_1013 = _decoder_T_607 ? 3'h4 : _decoder_T_1012; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_1014 = _decoder_T_605 ? 3'h2 : _decoder_T_1013; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_1015 = _decoder_T_603 ? 3'h2 : _decoder_T_1014; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_1016 = _decoder_T_601 ? 3'h4 : _decoder_T_1015; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_1017 = _decoder_T_599 ? 3'h4 : _decoder_T_1016; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_1018 = _decoder_T_597 ? 3'h4 : _decoder_T_1017; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_1019 = _decoder_T_595 ? 3'h4 : _decoder_T_1018; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_1020 = _decoder_T_593 ? 3'h2 : _decoder_T_1019; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_1021 = _decoder_T_591 ? 3'h1 : _decoder_T_1020; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_1022 = _decoder_T_589 ? 3'h2 : _decoder_T_1021; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_1023 = _decoder_T_587 ? 3'h1 : _decoder_T_1022; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_1024 = _decoder_T_585 ? 3'h2 : _decoder_T_1023; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_1025 = _decoder_T_583 ? 3'h2 : _decoder_T_1024; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_1026 = _decoder_T_581 ? 3'h2 : _decoder_T_1025; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_1027 = _decoder_T_579 ? 3'h1 : _decoder_T_1026; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_1028 = _decoder_T_577 ? 3'h2 : _decoder_T_1027; // @[Lookup.scala 33:37]
  wire [2:0] _decoder_T_1029 = _decoder_T_575 ? 3'h1 : _decoder_T_1028; // @[Lookup.scala 33:37]
  wire [2:0] decoder_5_1 = _decoder_T_573 ? 3'h2 : _decoder_T_1029; // @[Lookup.scala 33:37]
  wire  _decoder_T_1047 = _decoder_T_647 ? 1'h0 : _decoder_T_655 | (_decoder_T_657 | (_decoder_T_659 | (_decoder_T_661
     | (_decoder_T_663 | (_decoder_T_665 | _decoder_T_667))))); // @[Lookup.scala 33:37]
  wire  _decoder_T_1048 = _decoder_T_643 ? 1'h0 : _decoder_T_1047; // @[Lookup.scala 33:37]
  wire  _decoder_T_1049 = _decoder_T_649 ? 1'h0 : _decoder_T_1048; // @[Lookup.scala 33:37]
  wire  _decoder_T_1050 = _decoder_T_647 ? 1'h0 : _decoder_T_1049; // @[Lookup.scala 33:37]
  wire  _decoder_T_1051 = _decoder_T_645 ? 1'h0 : _decoder_T_1050; // @[Lookup.scala 33:37]
  wire  _decoder_T_1052 = _decoder_T_643 ? 1'h0 : _decoder_T_1051; // @[Lookup.scala 33:37]
  wire  _decoder_T_1053 = _decoder_T_641 ? 1'h0 : _decoder_T_1052; // @[Lookup.scala 33:37]
  wire  _decoder_T_1054 = _decoder_T_639 ? 1'h0 : _decoder_T_1053; // @[Lookup.scala 33:37]
  wire  _decoder_T_1055 = _decoder_T_637 ? 1'h0 : _decoder_T_1054; // @[Lookup.scala 33:37]
  wire  _decoder_T_1056 = _decoder_T_635 ? 1'h0 : _decoder_T_1055; // @[Lookup.scala 33:37]
  wire  _decoder_T_1057 = _decoder_T_633 ? 1'h0 : _decoder_T_1056; // @[Lookup.scala 33:37]
  wire  _decoder_T_1058 = _decoder_T_631 ? 1'h0 : _decoder_T_1057; // @[Lookup.scala 33:37]
  wire  _decoder_T_1059 = _decoder_T_629 ? 1'h0 : _decoder_T_1058; // @[Lookup.scala 33:37]
  wire  _decoder_T_1060 = _decoder_T_627 ? 1'h0 : _decoder_T_1059; // @[Lookup.scala 33:37]
  wire  _decoder_T_1061 = _decoder_T_625 ? 1'h0 : _decoder_T_1060; // @[Lookup.scala 33:37]
  wire  _decoder_T_1062 = _decoder_T_623 ? 1'h0 : _decoder_T_1061; // @[Lookup.scala 33:37]
  wire  _decoder_T_1063 = _decoder_T_621 ? 1'h0 : _decoder_T_1062; // @[Lookup.scala 33:37]
  wire  _decoder_T_1064 = _decoder_T_619 ? 1'h0 : _decoder_T_1063; // @[Lookup.scala 33:37]
  wire  _decoder_T_1065 = _decoder_T_617 ? 1'h0 : _decoder_T_1064; // @[Lookup.scala 33:37]
  wire  _decoder_T_1066 = _decoder_T_615 ? 1'h0 : _decoder_T_1065; // @[Lookup.scala 33:37]
  wire  _decoder_T_1067 = _decoder_T_613 ? 1'h0 : _decoder_T_1066; // @[Lookup.scala 33:37]
  wire  _decoder_T_1068 = _decoder_T_611 ? 1'h0 : _decoder_T_1067; // @[Lookup.scala 33:37]
  wire  _decoder_T_1069 = _decoder_T_609 ? 1'h0 : _decoder_T_1068; // @[Lookup.scala 33:37]
  wire  _decoder_T_1070 = _decoder_T_607 ? 1'h0 : _decoder_T_1069; // @[Lookup.scala 33:37]
  wire  _decoder_T_1071 = _decoder_T_605 ? 1'h0 : _decoder_T_1070; // @[Lookup.scala 33:37]
  wire  _decoder_T_1072 = _decoder_T_603 ? 1'h0 : _decoder_T_1071; // @[Lookup.scala 33:37]
  wire  _decoder_T_1073 = _decoder_T_601 ? 1'h0 : _decoder_T_1072; // @[Lookup.scala 33:37]
  wire  _decoder_T_1074 = _decoder_T_599 ? 1'h0 : _decoder_T_1073; // @[Lookup.scala 33:37]
  wire  _decoder_T_1075 = _decoder_T_597 ? 1'h0 : _decoder_T_1074; // @[Lookup.scala 33:37]
  wire  _decoder_T_1076 = _decoder_T_595 ? 1'h0 : _decoder_T_1075; // @[Lookup.scala 33:37]
  wire  _decoder_T_1077 = _decoder_T_593 ? 1'h0 : _decoder_T_1076; // @[Lookup.scala 33:37]
  wire  _decoder_T_1078 = _decoder_T_591 ? 1'h0 : _decoder_T_1077; // @[Lookup.scala 33:37]
  wire  _decoder_T_1079 = _decoder_T_589 ? 1'h0 : _decoder_T_1078; // @[Lookup.scala 33:37]
  wire  _decoder_T_1080 = _decoder_T_587 ? 1'h0 : _decoder_T_1079; // @[Lookup.scala 33:37]
  wire  _decoder_T_1081 = _decoder_T_585 ? 1'h0 : _decoder_T_1080; // @[Lookup.scala 33:37]
  wire  _decoder_T_1082 = _decoder_T_583 ? 1'h0 : _decoder_T_1081; // @[Lookup.scala 33:37]
  wire  _decoder_T_1083 = _decoder_T_581 ? 1'h0 : _decoder_T_1082; // @[Lookup.scala 33:37]
  wire  _decoder_T_1084 = _decoder_T_579 ? 1'h0 : _decoder_T_1083; // @[Lookup.scala 33:37]
  wire  _decoder_T_1085 = _decoder_T_577 ? 1'h0 : _decoder_T_1084; // @[Lookup.scala 33:37]
  wire [4:0] rs_1 = io_fb_inst_bank_bits_data_1_inst[25:21]; // @[Decode.scala 34:27]
  wire [4:0] rt_1 = io_fb_inst_bank_bits_data_1_inst[20:16]; // @[Decode.scala 35:27]
  wire [4:0] rd_1 = io_fb_inst_bank_bits_data_1_inst[15:11]; // @[Decode.scala 36:27]
  wire [15:0] rename_info_1_imm_data_lo = io_fb_inst_bank_bits_data_1_inst[15:0]; // @[Decode.scala 37:27]
  wire [25:0] rename_info_1_imm_data_lo_1 = io_fb_inst_bank_bits_data_1_inst[25:0]; // @[Decode.scala 38:27]
  wire [4:0] rename_info_1_imm_data_lo_2 = io_fb_inst_bank_bits_data_1_inst[10:6]; // @[Decode.scala 39:27]
  wire  rename_info_1_need_imm = decoder_2_1 != 3'h4; // @[Decode.scala 46:25]
  wire [4:0] _rename_info_1_op1_addr_T_6 = 3'h0 == decoder_3_1 ? rs_1 : 5'h0; // @[Mux.scala 80:57]
  wire [4:0] _rename_info_1_op1_addr_T_8 = 3'h1 == decoder_3_1 ? rt_1 : _rename_info_1_op1_addr_T_6; // @[Mux.scala 80:57]
  wire [4:0] _rename_info_1_op1_addr_T_10 = 3'h2 == decoder_3_1 ? rd_1 : _rename_info_1_op1_addr_T_8; // @[Mux.scala 80:57]
  wire [4:0] rename_info_1_op1_addr = 3'h3 == decoder_3_1 ? 5'h1f : _rename_info_1_op1_addr_T_10; // @[Mux.scala 80:57]
  wire [4:0] _rename_info_1_op2_addr_T_6 = 3'h0 == decoder_4_1 ? rs_1 : 5'h0; // @[Mux.scala 80:57]
  wire [4:0] _rename_info_1_op2_addr_T_8 = 3'h1 == decoder_4_1 ? rt_1 : _rename_info_1_op2_addr_T_6; // @[Mux.scala 80:57]
  wire [4:0] _rename_info_1_op2_addr_T_10 = 3'h2 == decoder_4_1 ? rd_1 : _rename_info_1_op2_addr_T_8; // @[Mux.scala 80:57]
  wire [4:0] rename_info_1_op2_addr = 3'h3 == decoder_4_1 ? 5'h1f : _rename_info_1_op2_addr_T_10; // @[Mux.scala 80:57]
  wire [4:0] _rename_info_1_des_addr_T_6 = 3'h0 == decoder_5_1 ? rs_1 : 5'h0; // @[Mux.scala 80:57]
  wire [4:0] _rename_info_1_des_addr_T_8 = 3'h1 == decoder_5_1 ? rt_1 : _rename_info_1_des_addr_T_6; // @[Mux.scala 80:57]
  wire [4:0] _rename_info_1_des_addr_T_10 = 3'h2 == decoder_5_1 ? rd_1 : _rename_info_1_des_addr_T_8; // @[Mux.scala 80:57]
  wire [4:0] rename_info_1_des_addr = 3'h3 == decoder_5_1 ? 5'h1f : _rename_info_1_des_addr_T_10; // @[Mux.scala 80:57]
  wire [15:0] rename_info_1_imm_data_hi = rename_info_1_imm_data_lo[15] ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _rename_info_1_imm_data_T_4 = {rename_info_1_imm_data_hi,rename_info_1_imm_data_lo}; // @[Cat.scala 30:58]
  wire [31:0] _rename_info_1_imm_data_T_6 = {16'h0,rename_info_1_imm_data_lo}; // @[Cat.scala 30:58]
  wire [31:0] _rename_info_1_imm_data_T_8 = {27'h0,rename_info_1_imm_data_lo_2}; // @[Cat.scala 30:58]
  wire [35:0] _rename_info_1_imm_data_T_10 = {10'h0,rename_info_1_imm_data_lo_1}; // @[Cat.scala 30:58]
  wire [31:0] _rename_info_1_imm_data_T_12 = 3'h1 == decoder_2_1 ? _rename_info_1_imm_data_T_4 : 32'h0; // @[Mux.scala 80:57]
  wire [31:0] _rename_info_1_imm_data_T_14 = 3'h0 == decoder_2_1 ? _rename_info_1_imm_data_T_6 :
    _rename_info_1_imm_data_T_12; // @[Mux.scala 80:57]
  wire [31:0] _rename_info_1_imm_data_T_16 = 3'h2 == decoder_2_1 ? _rename_info_1_imm_data_T_8 :
    _rename_info_1_imm_data_T_14; // @[Mux.scala 80:57]
  wire [35:0] _rename_info_1_imm_data_T_18 = 3'h3 == decoder_2_1 ? _rename_info_1_imm_data_T_10 : {{4'd0},
    _rename_info_1_imm_data_T_16}; // @[Mux.scala 80:57]
  reg [2:0] rob_allocate_info_bits_0_rob_idx; // @[Decode.scala 115:35]
  reg  rob_allocate_info_bits_0_inst_valid; // @[Decode.scala 115:35]
  reg [31:0] rob_allocate_info_bits_0_inst_addr; // @[Decode.scala 115:35]
  reg [5:0] rob_allocate_info_bits_0_uop; // @[Decode.scala 115:35]
  reg [2:0] rob_allocate_info_bits_0_unit_sel; // @[Decode.scala 115:35]
  reg  rob_allocate_info_bits_0_need_imm; // @[Decode.scala 115:35]
  reg [31:0] rob_allocate_info_bits_0_commit_addr; // @[Decode.scala 115:35]
  reg [3:0] rob_allocate_info_bits_0_gh_info; // @[Decode.scala 115:35]
  reg [31:0] rob_allocate_info_bits_0_imm_data; // @[Decode.scala 115:35]
  reg  rob_allocate_info_bits_0_flush_on_commit; // @[Decode.scala 115:35]
  reg  rob_allocate_info_bits_0_predict_taken; // @[Decode.scala 115:35]
  reg [2:0] rob_allocate_info_bits_1_rob_idx; // @[Decode.scala 115:35]
  reg  rob_allocate_info_bits_1_inst_valid; // @[Decode.scala 115:35]
  reg [31:0] rob_allocate_info_bits_1_inst_addr; // @[Decode.scala 115:35]
  reg [5:0] rob_allocate_info_bits_1_uop; // @[Decode.scala 115:35]
  reg [2:0] rob_allocate_info_bits_1_unit_sel; // @[Decode.scala 115:35]
  reg  rob_allocate_info_bits_1_need_imm; // @[Decode.scala 115:35]
  reg [31:0] rob_allocate_info_bits_1_commit_addr; // @[Decode.scala 115:35]
  reg [3:0] rob_allocate_info_bits_1_gh_info; // @[Decode.scala 115:35]
  reg [31:0] rob_allocate_info_bits_1_imm_data; // @[Decode.scala 115:35]
  reg  rob_allocate_info_bits_1_flush_on_commit; // @[Decode.scala 115:35]
  reg  rob_allocate_info_bits_1_predict_taken; // @[Decode.scala 115:35]
  reg  rob_allocate_info_valid; // @[Decode.scala 116:40]
  wire  _GEN_0 = io_need_flush ? 1'h0 : io_rob_allocate_allocate_resp_bits_enq_valid_mask_0; // @[Decode.scala 153:22 Decode.scala 82:14 Decode.scala 140:34]
  wire [4:0] _GEN_1 = io_need_flush ? 5'h0 : rename_info_0_op1_addr; // @[Decode.scala 153:22 Decode.scala 83:14 Decode.scala 141:34]
  wire [4:0] _GEN_2 = io_need_flush ? 5'h0 : rename_info_0_op2_addr; // @[Decode.scala 153:22 Decode.scala 84:14 Decode.scala 142:34]
  wire [4:0] _GEN_3 = io_need_flush ? 5'h0 : rename_info_0_des_addr; // @[Decode.scala 153:22 Decode.scala 85:14 Decode.scala 143:34]
  wire [2:0] _GEN_4 = io_need_flush ? 3'h0 : io_rob_allocate_allocate_resp_bits_rob_idx_0; // @[Decode.scala 153:22 Decode.scala 86:14 Decode.scala 144:34]
  wire  _GEN_5 = io_need_flush ? 1'h0 : io_rob_allocate_allocate_resp_bits_enq_valid_mask_1; // @[Decode.scala 153:22 Decode.scala 82:14 Decode.scala 140:34]
  wire [4:0] _GEN_6 = io_need_flush ? 5'h0 : rename_info_1_op1_addr; // @[Decode.scala 153:22 Decode.scala 83:14 Decode.scala 141:34]
  wire [4:0] _GEN_7 = io_need_flush ? 5'h0 : rename_info_1_op2_addr; // @[Decode.scala 153:22 Decode.scala 84:14 Decode.scala 142:34]
  wire [4:0] _GEN_8 = io_need_flush ? 5'h0 : rename_info_1_des_addr; // @[Decode.scala 153:22 Decode.scala 85:14 Decode.scala 143:34]
  wire [2:0] _GEN_9 = io_need_flush ? 3'h0 : io_rob_allocate_allocate_resp_bits_rob_idx_1; // @[Decode.scala 153:22 Decode.scala 86:14 Decode.scala 144:34]
  wire [31:0] rename_info_0_imm_data = _rename_info_0_imm_data_T_18[31:0]; // @[Decode.scala 105:25 Decode.scala 65:14]
  wire [31:0] rename_info_1_imm_data = _rename_info_1_imm_data_T_18[31:0]; // @[Decode.scala 105:25 Decode.scala 65:14]
  assign io_fb_resp_deq_valid_0 = io_rob_allocate_allocate_resp_bits_enq_valid_mask_0; // @[Decode.scala 151:23]
  assign io_fb_resp_deq_valid_1 = io_rob_allocate_allocate_resp_bits_enq_valid_mask_1; // @[Decode.scala 151:23]
  assign io_rob_allocate_allocate_req_valid = io_fb_inst_bank_valid; // @[Decode.scala 113:37]
  assign io_rob_allocate_allocate_req_bits_0 = io_fb_inst_bank_bits_data_0_is_valid; // @[Decode.scala 112:46 Decode.scala 112:46]
  assign io_rob_allocate_allocate_req_bits_1 = io_fb_inst_bank_bits_data_1_is_valid; // @[Decode.scala 112:46 Decode.scala 112:46]
  assign io_rob_allocate_allocate_info_valid = rob_allocate_info_valid; // @[Decode.scala 120:38]
  assign io_rob_allocate_allocate_info_bits_0_rob_idx = rob_allocate_info_bits_0_rob_idx; // @[Decode.scala 119:37]
  assign io_rob_allocate_allocate_info_bits_0_inst_valid = rob_allocate_info_bits_0_inst_valid; // @[Decode.scala 119:37]
  assign io_rob_allocate_allocate_info_bits_0_inst_addr = rob_allocate_info_bits_0_inst_addr; // @[Decode.scala 119:37]
  assign io_rob_allocate_allocate_info_bits_0_uop = rob_allocate_info_bits_0_uop; // @[Decode.scala 119:37]
  assign io_rob_allocate_allocate_info_bits_0_unit_sel = rob_allocate_info_bits_0_unit_sel; // @[Decode.scala 119:37]
  assign io_rob_allocate_allocate_info_bits_0_need_imm = rob_allocate_info_bits_0_need_imm; // @[Decode.scala 119:37]
  assign io_rob_allocate_allocate_info_bits_0_commit_addr = rob_allocate_info_bits_0_commit_addr; // @[Decode.scala 119:37]
  assign io_rob_allocate_allocate_info_bits_0_gh_info = rob_allocate_info_bits_0_gh_info; // @[Decode.scala 119:37]
  assign io_rob_allocate_allocate_info_bits_0_imm_data = rob_allocate_info_bits_0_imm_data; // @[Decode.scala 119:37]
  assign io_rob_allocate_allocate_info_bits_0_flush_on_commit = rob_allocate_info_bits_0_flush_on_commit; // @[Decode.scala 119:37]
  assign io_rob_allocate_allocate_info_bits_0_predict_taken = rob_allocate_info_bits_0_predict_taken; // @[Decode.scala 119:37]
  assign io_rob_allocate_allocate_info_bits_1_rob_idx = rob_allocate_info_bits_1_rob_idx; // @[Decode.scala 119:37]
  assign io_rob_allocate_allocate_info_bits_1_inst_valid = rob_allocate_info_bits_1_inst_valid; // @[Decode.scala 119:37]
  assign io_rob_allocate_allocate_info_bits_1_inst_addr = rob_allocate_info_bits_1_inst_addr; // @[Decode.scala 119:37]
  assign io_rob_allocate_allocate_info_bits_1_uop = rob_allocate_info_bits_1_uop; // @[Decode.scala 119:37]
  assign io_rob_allocate_allocate_info_bits_1_unit_sel = rob_allocate_info_bits_1_unit_sel; // @[Decode.scala 119:37]
  assign io_rob_allocate_allocate_info_bits_1_need_imm = rob_allocate_info_bits_1_need_imm; // @[Decode.scala 119:37]
  assign io_rob_allocate_allocate_info_bits_1_commit_addr = rob_allocate_info_bits_1_commit_addr; // @[Decode.scala 119:37]
  assign io_rob_allocate_allocate_info_bits_1_gh_info = rob_allocate_info_bits_1_gh_info; // @[Decode.scala 119:37]
  assign io_rob_allocate_allocate_info_bits_1_imm_data = rob_allocate_info_bits_1_imm_data; // @[Decode.scala 119:37]
  assign io_rob_allocate_allocate_info_bits_1_flush_on_commit = rob_allocate_info_bits_1_flush_on_commit; // @[Decode.scala 119:37]
  assign io_rob_allocate_allocate_info_bits_1_predict_taken = rob_allocate_info_bits_1_predict_taken; // @[Decode.scala 119:37]
  assign io_rename_info_valid = io_need_flush ? 1'h0 : io_fb_inst_bank_valid & io_rob_allocate_allocate_resp_valid; // @[Decode.scala 153:22 Decode.scala 155:22 Decode.scala 146:21]
  assign io_rename_info_bits_0_is_valid = reset ? 1'h0 : _GEN_0; // @[Decode.scala 160:23 Decode.scala 82:14]
  assign io_rename_info_bits_0_op1_addr = reset ? 5'h0 : _GEN_1; // @[Decode.scala 160:23 Decode.scala 83:14]
  assign io_rename_info_bits_0_op2_addr = reset ? 5'h0 : _GEN_2; // @[Decode.scala 160:23 Decode.scala 84:14]
  assign io_rename_info_bits_0_des_addr = reset ? 5'h0 : _GEN_3; // @[Decode.scala 160:23 Decode.scala 85:14]
  assign io_rename_info_bits_0_des_rob = reset ? 3'h0 : _GEN_4; // @[Decode.scala 160:23 Decode.scala 86:14]
  assign io_rename_info_bits_1_is_valid = reset ? 1'h0 : _GEN_5; // @[Decode.scala 160:23 Decode.scala 82:14]
  assign io_rename_info_bits_1_op1_addr = reset ? 5'h0 : _GEN_6; // @[Decode.scala 160:23 Decode.scala 83:14]
  assign io_rename_info_bits_1_op2_addr = reset ? 5'h0 : _GEN_7; // @[Decode.scala 160:23 Decode.scala 84:14]
  assign io_rename_info_bits_1_des_addr = reset ? 5'h0 : _GEN_8; // @[Decode.scala 160:23 Decode.scala 85:14]
  assign io_rename_info_bits_1_des_rob = reset ? 3'h0 : _GEN_9; // @[Decode.scala 160:23 Decode.scala 86:14]
  always @(posedge clock) begin
    if (reset) begin // @[Decode.scala 160:23]
      rob_allocate_info_bits_0_rob_idx <= 3'h0; // @[Decode.scala 86:14]
    end else if (io_need_flush) begin // @[Decode.scala 153:22]
      rob_allocate_info_bits_0_rob_idx <= 3'h0; // @[Decode.scala 86:14]
    end else begin
      rob_allocate_info_bits_0_rob_idx <= io_rob_allocate_allocate_resp_bits_rob_idx_0; // @[Decode.scala 144:34]
    end
    if (reset) begin // @[Decode.scala 160:23]
      rob_allocate_info_bits_0_inst_valid <= 1'h0; // @[Decode.scala 82:14]
    end else if (io_need_flush) begin // @[Decode.scala 153:22]
      rob_allocate_info_bits_0_inst_valid <= 1'h0; // @[Decode.scala 82:14]
    end else begin
      rob_allocate_info_bits_0_inst_valid <= io_rob_allocate_allocate_resp_bits_enq_valid_mask_0; // @[Decode.scala 140:34]
    end
    if (reset) begin // @[Decode.scala 160:23]
      rob_allocate_info_bits_0_inst_addr <= 32'h0; // @[Rob.scala 90:21]
    end else if (io_need_flush) begin // @[Decode.scala 153:22]
      rob_allocate_info_bits_0_inst_addr <= 32'h0; // @[Rob.scala 90:21]
    end else begin
      rob_allocate_info_bits_0_inst_addr <= io_fb_inst_bank_bits_data_0_inst_addr; // @[Decode.scala 125:41]
    end
    if (reset) begin // @[Decode.scala 160:23]
      rob_allocate_info_bits_0_uop <= 6'h0; // @[Rob.scala 91:21]
    end else if (io_need_flush) begin // @[Decode.scala 153:22]
      rob_allocate_info_bits_0_uop <= 6'h0; // @[Rob.scala 91:21]
    end else if (_decoder_T_1) begin // @[Lookup.scala 33:37]
      rob_allocate_info_bits_0_uop <= 6'h1;
    end else if (_decoder_T_3) begin // @[Lookup.scala 33:37]
      rob_allocate_info_bits_0_uop <= 6'h1;
    end else begin
      rob_allocate_info_bits_0_uop <= _decoder_T_171;
    end
    if (reset) begin // @[Decode.scala 160:23]
      rob_allocate_info_bits_0_unit_sel <= 3'h0; // @[Rob.scala 92:21]
    end else if (io_need_flush) begin // @[Decode.scala 153:22]
      rob_allocate_info_bits_0_unit_sel <= 3'h0; // @[Rob.scala 92:21]
    end else if (_decoder_T_1) begin // @[Lookup.scala 33:37]
      rob_allocate_info_bits_0_unit_sel <= 3'h1;
    end else if (_decoder_T_3) begin // @[Lookup.scala 33:37]
      rob_allocate_info_bits_0_unit_sel <= 3'h1;
    end else begin
      rob_allocate_info_bits_0_unit_sel <= _decoder_T_228;
    end
    if (reset) begin // @[Decode.scala 160:23]
      rob_allocate_info_bits_0_need_imm <= 1'h0; // @[Rob.scala 93:21]
    end else if (io_need_flush) begin // @[Decode.scala 153:22]
      rob_allocate_info_bits_0_need_imm <= 1'h0; // @[Rob.scala 93:21]
    end else begin
      rob_allocate_info_bits_0_need_imm <= rename_info_0_need_imm; // @[Decode.scala 137:40]
    end
    if (reset) begin // @[Decode.scala 160:23]
      rob_allocate_info_bits_0_commit_addr <= 32'h0; // @[Rob.scala 94:21]
    end else if (io_need_flush) begin // @[Decode.scala 153:22]
      rob_allocate_info_bits_0_commit_addr <= 32'h0; // @[Rob.scala 94:21]
    end else begin
      rob_allocate_info_bits_0_commit_addr <= {{27'd0}, rename_info_0_des_addr}; // @[Decode.scala 126:43]
    end
    if (reset) begin // @[Decode.scala 160:23]
      rob_allocate_info_bits_0_gh_info <= 4'h0; // @[Rob.scala 99:21]
    end else if (io_need_flush) begin // @[Decode.scala 153:22]
      rob_allocate_info_bits_0_gh_info <= 4'h0; // @[Rob.scala 99:21]
    end else begin
      rob_allocate_info_bits_0_gh_info <= io_fb_inst_bank_bits_data_0_gh_backup; // @[Decode.scala 132:39]
    end
    if (reset) begin // @[Decode.scala 160:23]
      rob_allocate_info_bits_0_imm_data <= 32'h0; // @[Rob.scala 100:21]
    end else if (io_need_flush) begin // @[Decode.scala 153:22]
      rob_allocate_info_bits_0_imm_data <= 32'h0; // @[Rob.scala 100:21]
    end else begin
      rob_allocate_info_bits_0_imm_data <= rename_info_0_imm_data; // @[Decode.scala 133:40]
    end
    if (reset) begin // @[Decode.scala 160:23]
      rob_allocate_info_bits_0_flush_on_commit <= 1'h0; // @[Rob.scala 101:21]
    end else if (io_need_flush) begin // @[Decode.scala 153:22]
      rob_allocate_info_bits_0_flush_on_commit <= 1'h0; // @[Rob.scala 101:21]
    end else if (_decoder_T_1) begin // @[Lookup.scala 33:37]
      rob_allocate_info_bits_0_flush_on_commit <= 1'h0;
    end else if (_decoder_T_3) begin // @[Lookup.scala 33:37]
      rob_allocate_info_bits_0_flush_on_commit <= 1'h0;
    end else begin
      rob_allocate_info_bits_0_flush_on_commit <= _decoder_T_513;
    end
    if (reset) begin // @[Decode.scala 160:23]
      rob_allocate_info_bits_0_predict_taken <= 1'h0; // @[Rob.scala 102:21]
    end else if (io_need_flush) begin // @[Decode.scala 153:22]
      rob_allocate_info_bits_0_predict_taken <= 1'h0; // @[Rob.scala 102:21]
    end else begin
      rob_allocate_info_bits_0_predict_taken <= io_fb_inst_bank_bits_data_0_predict_taken; // @[Decode.scala 131:45]
    end
    if (reset) begin // @[Decode.scala 160:23]
      rob_allocate_info_bits_1_rob_idx <= 3'h0; // @[Decode.scala 86:14]
    end else if (io_need_flush) begin // @[Decode.scala 153:22]
      rob_allocate_info_bits_1_rob_idx <= 3'h0; // @[Decode.scala 86:14]
    end else begin
      rob_allocate_info_bits_1_rob_idx <= io_rob_allocate_allocate_resp_bits_rob_idx_1; // @[Decode.scala 144:34]
    end
    if (reset) begin // @[Decode.scala 160:23]
      rob_allocate_info_bits_1_inst_valid <= 1'h0; // @[Decode.scala 82:14]
    end else if (io_need_flush) begin // @[Decode.scala 153:22]
      rob_allocate_info_bits_1_inst_valid <= 1'h0; // @[Decode.scala 82:14]
    end else begin
      rob_allocate_info_bits_1_inst_valid <= io_rob_allocate_allocate_resp_bits_enq_valid_mask_1; // @[Decode.scala 140:34]
    end
    if (reset) begin // @[Decode.scala 160:23]
      rob_allocate_info_bits_1_inst_addr <= 32'h0; // @[Rob.scala 90:21]
    end else if (io_need_flush) begin // @[Decode.scala 153:22]
      rob_allocate_info_bits_1_inst_addr <= 32'h0; // @[Rob.scala 90:21]
    end else begin
      rob_allocate_info_bits_1_inst_addr <= io_fb_inst_bank_bits_data_1_inst_addr; // @[Decode.scala 125:41]
    end
    if (reset) begin // @[Decode.scala 160:23]
      rob_allocate_info_bits_1_uop <= 6'h0; // @[Rob.scala 91:21]
    end else if (io_need_flush) begin // @[Decode.scala 153:22]
      rob_allocate_info_bits_1_uop <= 6'h0; // @[Rob.scala 91:21]
    end else if (_decoder_T_573) begin // @[Lookup.scala 33:37]
      rob_allocate_info_bits_1_uop <= 6'h1;
    end else if (_decoder_T_575) begin // @[Lookup.scala 33:37]
      rob_allocate_info_bits_1_uop <= 6'h1;
    end else begin
      rob_allocate_info_bits_1_uop <= _decoder_T_743;
    end
    if (reset) begin // @[Decode.scala 160:23]
      rob_allocate_info_bits_1_unit_sel <= 3'h0; // @[Rob.scala 92:21]
    end else if (io_need_flush) begin // @[Decode.scala 153:22]
      rob_allocate_info_bits_1_unit_sel <= 3'h0; // @[Rob.scala 92:21]
    end else if (_decoder_T_573) begin // @[Lookup.scala 33:37]
      rob_allocate_info_bits_1_unit_sel <= 3'h1;
    end else if (_decoder_T_575) begin // @[Lookup.scala 33:37]
      rob_allocate_info_bits_1_unit_sel <= 3'h1;
    end else begin
      rob_allocate_info_bits_1_unit_sel <= _decoder_T_800;
    end
    if (reset) begin // @[Decode.scala 160:23]
      rob_allocate_info_bits_1_need_imm <= 1'h0; // @[Rob.scala 93:21]
    end else if (io_need_flush) begin // @[Decode.scala 153:22]
      rob_allocate_info_bits_1_need_imm <= 1'h0; // @[Rob.scala 93:21]
    end else begin
      rob_allocate_info_bits_1_need_imm <= rename_info_1_need_imm; // @[Decode.scala 137:40]
    end
    if (reset) begin // @[Decode.scala 160:23]
      rob_allocate_info_bits_1_commit_addr <= 32'h0; // @[Rob.scala 94:21]
    end else if (io_need_flush) begin // @[Decode.scala 153:22]
      rob_allocate_info_bits_1_commit_addr <= 32'h0; // @[Rob.scala 94:21]
    end else begin
      rob_allocate_info_bits_1_commit_addr <= {{27'd0}, rename_info_1_des_addr}; // @[Decode.scala 126:43]
    end
    if (reset) begin // @[Decode.scala 160:23]
      rob_allocate_info_bits_1_gh_info <= 4'h0; // @[Rob.scala 99:21]
    end else if (io_need_flush) begin // @[Decode.scala 153:22]
      rob_allocate_info_bits_1_gh_info <= 4'h0; // @[Rob.scala 99:21]
    end else begin
      rob_allocate_info_bits_1_gh_info <= io_fb_inst_bank_bits_data_1_gh_backup; // @[Decode.scala 132:39]
    end
    if (reset) begin // @[Decode.scala 160:23]
      rob_allocate_info_bits_1_imm_data <= 32'h0; // @[Rob.scala 100:21]
    end else if (io_need_flush) begin // @[Decode.scala 153:22]
      rob_allocate_info_bits_1_imm_data <= 32'h0; // @[Rob.scala 100:21]
    end else begin
      rob_allocate_info_bits_1_imm_data <= rename_info_1_imm_data; // @[Decode.scala 133:40]
    end
    if (reset) begin // @[Decode.scala 160:23]
      rob_allocate_info_bits_1_flush_on_commit <= 1'h0; // @[Rob.scala 101:21]
    end else if (io_need_flush) begin // @[Decode.scala 153:22]
      rob_allocate_info_bits_1_flush_on_commit <= 1'h0; // @[Rob.scala 101:21]
    end else if (_decoder_T_573) begin // @[Lookup.scala 33:37]
      rob_allocate_info_bits_1_flush_on_commit <= 1'h0;
    end else if (_decoder_T_575) begin // @[Lookup.scala 33:37]
      rob_allocate_info_bits_1_flush_on_commit <= 1'h0;
    end else begin
      rob_allocate_info_bits_1_flush_on_commit <= _decoder_T_1085;
    end
    if (reset) begin // @[Decode.scala 160:23]
      rob_allocate_info_bits_1_predict_taken <= 1'h0; // @[Rob.scala 102:21]
    end else if (io_need_flush) begin // @[Decode.scala 153:22]
      rob_allocate_info_bits_1_predict_taken <= 1'h0; // @[Rob.scala 102:21]
    end else begin
      rob_allocate_info_bits_1_predict_taken <= io_fb_inst_bank_bits_data_1_predict_taken; // @[Decode.scala 131:45]
    end
    if (reset) begin // @[Decode.scala 116:40]
      rob_allocate_info_valid <= 1'h0; // @[Decode.scala 116:40]
    end else if (io_need_flush) begin // @[Decode.scala 153:22]
      rob_allocate_info_valid <= 1'h0; // @[Decode.scala 157:28]
    end else begin
      rob_allocate_info_valid <= io_fb_inst_bank_valid; // @[Decode.scala 117:27]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  rob_allocate_info_bits_0_rob_idx = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  rob_allocate_info_bits_0_inst_valid = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  rob_allocate_info_bits_0_inst_addr = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  rob_allocate_info_bits_0_uop = _RAND_3[5:0];
  _RAND_4 = {1{`RANDOM}};
  rob_allocate_info_bits_0_unit_sel = _RAND_4[2:0];
  _RAND_5 = {1{`RANDOM}};
  rob_allocate_info_bits_0_need_imm = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  rob_allocate_info_bits_0_commit_addr = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  rob_allocate_info_bits_0_gh_info = _RAND_7[3:0];
  _RAND_8 = {1{`RANDOM}};
  rob_allocate_info_bits_0_imm_data = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  rob_allocate_info_bits_0_flush_on_commit = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  rob_allocate_info_bits_0_predict_taken = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  rob_allocate_info_bits_1_rob_idx = _RAND_11[2:0];
  _RAND_12 = {1{`RANDOM}};
  rob_allocate_info_bits_1_inst_valid = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  rob_allocate_info_bits_1_inst_addr = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  rob_allocate_info_bits_1_uop = _RAND_14[5:0];
  _RAND_15 = {1{`RANDOM}};
  rob_allocate_info_bits_1_unit_sel = _RAND_15[2:0];
  _RAND_16 = {1{`RANDOM}};
  rob_allocate_info_bits_1_need_imm = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  rob_allocate_info_bits_1_commit_addr = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  rob_allocate_info_bits_1_gh_info = _RAND_18[3:0];
  _RAND_19 = {1{`RANDOM}};
  rob_allocate_info_bits_1_imm_data = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  rob_allocate_info_bits_1_flush_on_commit = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  rob_allocate_info_bits_1_predict_taken = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  rob_allocate_info_valid = _RAND_22[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Rename(
  input         clock,
  input         reset,
  input         io_rename_info_valid,
  input         io_rename_info_bits_0_is_valid,
  input  [4:0]  io_rename_info_bits_0_op1_addr,
  input  [4:0]  io_rename_info_bits_0_op2_addr,
  input  [4:0]  io_rename_info_bits_0_des_addr,
  input  [2:0]  io_rename_info_bits_0_des_rob,
  input         io_rename_info_bits_1_is_valid,
  input  [4:0]  io_rename_info_bits_1_op1_addr,
  input  [4:0]  io_rename_info_bits_1_op2_addr,
  input  [4:0]  io_rename_info_bits_1_des_addr,
  input  [2:0]  io_rename_info_bits_1_des_rob,
  input         io_rob_commit_0_valid,
  input  [2:0]  io_rob_commit_0_bits_des_rob,
  input  [4:0]  io_rob_commit_0_bits_commit_addr,
  input         io_rob_commit_1_valid,
  input  [2:0]  io_rob_commit_1_bits_des_rob,
  input  [4:0]  io_rob_commit_1_bits_commit_addr,
  output [4:0]  io_reg_read_0_op1_addr,
  output [4:0]  io_reg_read_0_op2_addr,
  input  [31:0] io_reg_read_0_op1_data,
  input  [31:0] io_reg_read_0_op2_data,
  output [4:0]  io_reg_read_1_op1_addr,
  output [4:0]  io_reg_read_1_op2_addr,
  input  [31:0] io_reg_read_1_op1_data,
  input  [31:0] io_reg_read_1_op2_data,
  output        io_rob_init_info_valid,
  output        io_rob_init_info_bits_0_is_valid,
  output [2:0]  io_rob_init_info_bits_0_des_rob,
  output [2:0]  io_rob_init_info_bits_0_op1_rob,
  output [2:0]  io_rob_init_info_bits_0_op2_rob,
  output [31:0] io_rob_init_info_bits_0_op1_regData,
  output [31:0] io_rob_init_info_bits_0_op2_regData,
  output        io_rob_init_info_bits_0_op1_in_rob,
  output        io_rob_init_info_bits_0_op2_in_rob,
  output        io_rob_init_info_bits_1_is_valid,
  output [2:0]  io_rob_init_info_bits_1_des_rob,
  output [2:0]  io_rob_init_info_bits_1_op1_rob,
  output [2:0]  io_rob_init_info_bits_1_op2_rob,
  output [31:0] io_rob_init_info_bits_1_op1_regData,
  output [31:0] io_rob_init_info_bits_1_op2_regData,
  output        io_rob_init_info_bits_1_op1_in_rob,
  output        io_rob_init_info_bits_1_op2_in_rob,
  input         io_need_flush
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] busy_table; // @[Rename.scala 60:27]
  reg [2:0] map_table_1; // @[Rename.scala 61:26]
  reg [2:0] map_table_2; // @[Rename.scala 61:26]
  reg [2:0] map_table_3; // @[Rename.scala 61:26]
  reg [2:0] map_table_4; // @[Rename.scala 61:26]
  reg [2:0] map_table_5; // @[Rename.scala 61:26]
  reg [2:0] map_table_6; // @[Rename.scala 61:26]
  reg [2:0] map_table_7; // @[Rename.scala 61:26]
  reg [2:0] map_table_8; // @[Rename.scala 61:26]
  reg [2:0] map_table_9; // @[Rename.scala 61:26]
  reg [2:0] map_table_10; // @[Rename.scala 61:26]
  reg [2:0] map_table_11; // @[Rename.scala 61:26]
  reg [2:0] map_table_12; // @[Rename.scala 61:26]
  reg [2:0] map_table_13; // @[Rename.scala 61:26]
  reg [2:0] map_table_14; // @[Rename.scala 61:26]
  reg [2:0] map_table_15; // @[Rename.scala 61:26]
  reg [2:0] map_table_16; // @[Rename.scala 61:26]
  reg [2:0] map_table_17; // @[Rename.scala 61:26]
  reg [2:0] map_table_18; // @[Rename.scala 61:26]
  reg [2:0] map_table_19; // @[Rename.scala 61:26]
  reg [2:0] map_table_20; // @[Rename.scala 61:26]
  reg [2:0] map_table_21; // @[Rename.scala 61:26]
  reg [2:0] map_table_22; // @[Rename.scala 61:26]
  reg [2:0] map_table_23; // @[Rename.scala 61:26]
  reg [2:0] map_table_24; // @[Rename.scala 61:26]
  reg [2:0] map_table_25; // @[Rename.scala 61:26]
  reg [2:0] map_table_26; // @[Rename.scala 61:26]
  reg [2:0] map_table_27; // @[Rename.scala 61:26]
  reg [2:0] map_table_28; // @[Rename.scala 61:26]
  reg [2:0] map_table_29; // @[Rename.scala 61:26]
  reg [2:0] map_table_30; // @[Rename.scala 61:26]
  reg [2:0] map_table_31; // @[Rename.scala 61:26]
  wire [31:0] _will_busy_T = 32'h1 << io_rename_info_bits_0_des_addr; // @[OneHot.scala 58:35]
  wire  _will_busy_T_1 = io_rename_info_valid & io_rename_info_bits_0_is_valid; // @[Rename.scala 63:95]
  wire [31:0] _will_busy_T_3 = _will_busy_T_1 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _will_busy_T_4 = _will_busy_T & _will_busy_T_3; // @[Rename.scala 63:66]
  wire [31:0] _will_busy_T_5 = 32'h1 << io_rename_info_bits_1_des_addr; // @[OneHot.scala 58:35]
  wire  _will_busy_T_6 = io_rename_info_valid & io_rename_info_bits_1_is_valid; // @[Rename.scala 63:95]
  wire [31:0] _will_busy_T_8 = _will_busy_T_6 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _will_busy_T_9 = _will_busy_T_5 & _will_busy_T_8; // @[Rename.scala 63:66]
  wire [31:0] _will_busy_T_10 = _will_busy_T_4 | _will_busy_T_9; // @[Rename.scala 63:118]
  wire [31:0] will_busy = _will_busy_T_10 & 32'hfffffffe; // @[Rename.scala 63:121]
  wire [31:0] _busy_table_wb_T = 32'h1 << io_rob_commit_0_bits_commit_addr; // @[OneHot.scala 58:35]
  wire [2:0] _GEN_1 = 5'h1 == io_rob_commit_0_bits_commit_addr ? map_table_1 : 3'h0; // @[Rename.scala 64:117 Rename.scala 64:117]
  wire [2:0] _GEN_2 = 5'h2 == io_rob_commit_0_bits_commit_addr ? map_table_2 : _GEN_1; // @[Rename.scala 64:117 Rename.scala 64:117]
  wire [2:0] _GEN_3 = 5'h3 == io_rob_commit_0_bits_commit_addr ? map_table_3 : _GEN_2; // @[Rename.scala 64:117 Rename.scala 64:117]
  wire [2:0] _GEN_4 = 5'h4 == io_rob_commit_0_bits_commit_addr ? map_table_4 : _GEN_3; // @[Rename.scala 64:117 Rename.scala 64:117]
  wire [2:0] _GEN_5 = 5'h5 == io_rob_commit_0_bits_commit_addr ? map_table_5 : _GEN_4; // @[Rename.scala 64:117 Rename.scala 64:117]
  wire [2:0] _GEN_6 = 5'h6 == io_rob_commit_0_bits_commit_addr ? map_table_6 : _GEN_5; // @[Rename.scala 64:117 Rename.scala 64:117]
  wire [2:0] _GEN_7 = 5'h7 == io_rob_commit_0_bits_commit_addr ? map_table_7 : _GEN_6; // @[Rename.scala 64:117 Rename.scala 64:117]
  wire [2:0] _GEN_8 = 5'h8 == io_rob_commit_0_bits_commit_addr ? map_table_8 : _GEN_7; // @[Rename.scala 64:117 Rename.scala 64:117]
  wire [2:0] _GEN_9 = 5'h9 == io_rob_commit_0_bits_commit_addr ? map_table_9 : _GEN_8; // @[Rename.scala 64:117 Rename.scala 64:117]
  wire [2:0] _GEN_10 = 5'ha == io_rob_commit_0_bits_commit_addr ? map_table_10 : _GEN_9; // @[Rename.scala 64:117 Rename.scala 64:117]
  wire [2:0] _GEN_11 = 5'hb == io_rob_commit_0_bits_commit_addr ? map_table_11 : _GEN_10; // @[Rename.scala 64:117 Rename.scala 64:117]
  wire [2:0] _GEN_12 = 5'hc == io_rob_commit_0_bits_commit_addr ? map_table_12 : _GEN_11; // @[Rename.scala 64:117 Rename.scala 64:117]
  wire [2:0] _GEN_13 = 5'hd == io_rob_commit_0_bits_commit_addr ? map_table_13 : _GEN_12; // @[Rename.scala 64:117 Rename.scala 64:117]
  wire [2:0] _GEN_14 = 5'he == io_rob_commit_0_bits_commit_addr ? map_table_14 : _GEN_13; // @[Rename.scala 64:117 Rename.scala 64:117]
  wire [2:0] _GEN_15 = 5'hf == io_rob_commit_0_bits_commit_addr ? map_table_15 : _GEN_14; // @[Rename.scala 64:117 Rename.scala 64:117]
  wire [2:0] _GEN_16 = 5'h10 == io_rob_commit_0_bits_commit_addr ? map_table_16 : _GEN_15; // @[Rename.scala 64:117 Rename.scala 64:117]
  wire [2:0] _GEN_17 = 5'h11 == io_rob_commit_0_bits_commit_addr ? map_table_17 : _GEN_16; // @[Rename.scala 64:117 Rename.scala 64:117]
  wire [2:0] _GEN_18 = 5'h12 == io_rob_commit_0_bits_commit_addr ? map_table_18 : _GEN_17; // @[Rename.scala 64:117 Rename.scala 64:117]
  wire [2:0] _GEN_19 = 5'h13 == io_rob_commit_0_bits_commit_addr ? map_table_19 : _GEN_18; // @[Rename.scala 64:117 Rename.scala 64:117]
  wire [2:0] _GEN_20 = 5'h14 == io_rob_commit_0_bits_commit_addr ? map_table_20 : _GEN_19; // @[Rename.scala 64:117 Rename.scala 64:117]
  wire [2:0] _GEN_21 = 5'h15 == io_rob_commit_0_bits_commit_addr ? map_table_21 : _GEN_20; // @[Rename.scala 64:117 Rename.scala 64:117]
  wire [2:0] _GEN_22 = 5'h16 == io_rob_commit_0_bits_commit_addr ? map_table_22 : _GEN_21; // @[Rename.scala 64:117 Rename.scala 64:117]
  wire [2:0] _GEN_23 = 5'h17 == io_rob_commit_0_bits_commit_addr ? map_table_23 : _GEN_22; // @[Rename.scala 64:117 Rename.scala 64:117]
  wire [2:0] _GEN_24 = 5'h18 == io_rob_commit_0_bits_commit_addr ? map_table_24 : _GEN_23; // @[Rename.scala 64:117 Rename.scala 64:117]
  wire [2:0] _GEN_25 = 5'h19 == io_rob_commit_0_bits_commit_addr ? map_table_25 : _GEN_24; // @[Rename.scala 64:117 Rename.scala 64:117]
  wire [2:0] _GEN_26 = 5'h1a == io_rob_commit_0_bits_commit_addr ? map_table_26 : _GEN_25; // @[Rename.scala 64:117 Rename.scala 64:117]
  wire [2:0] _GEN_27 = 5'h1b == io_rob_commit_0_bits_commit_addr ? map_table_27 : _GEN_26; // @[Rename.scala 64:117 Rename.scala 64:117]
  wire [2:0] _GEN_28 = 5'h1c == io_rob_commit_0_bits_commit_addr ? map_table_28 : _GEN_27; // @[Rename.scala 64:117 Rename.scala 64:117]
  wire [2:0] _GEN_29 = 5'h1d == io_rob_commit_0_bits_commit_addr ? map_table_29 : _GEN_28; // @[Rename.scala 64:117 Rename.scala 64:117]
  wire [2:0] _GEN_30 = 5'h1e == io_rob_commit_0_bits_commit_addr ? map_table_30 : _GEN_29; // @[Rename.scala 64:117 Rename.scala 64:117]
  wire [2:0] _GEN_31 = 5'h1f == io_rob_commit_0_bits_commit_addr ? map_table_31 : _GEN_30; // @[Rename.scala 64:117 Rename.scala 64:117]
  wire  _busy_table_wb_T_2 = io_rob_commit_0_valid & io_rob_commit_0_bits_des_rob == _GEN_31; // @[Rename.scala 64:101]
  wire [31:0] _busy_table_wb_T_4 = _busy_table_wb_T_2 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _busy_table_wb_T_5 = _busy_table_wb_T & _busy_table_wb_T_4; // @[Rename.scala 64:85]
  wire [31:0] _busy_table_wb_T_6 = 32'h1 << io_rob_commit_1_bits_commit_addr; // @[OneHot.scala 58:35]
  wire [2:0] _GEN_33 = 5'h1 == io_rob_commit_1_bits_commit_addr ? map_table_1 : 3'h0; // @[Rename.scala 64:117 Rename.scala 64:117]
  wire [2:0] _GEN_34 = 5'h2 == io_rob_commit_1_bits_commit_addr ? map_table_2 : _GEN_33; // @[Rename.scala 64:117 Rename.scala 64:117]
  wire [2:0] _GEN_35 = 5'h3 == io_rob_commit_1_bits_commit_addr ? map_table_3 : _GEN_34; // @[Rename.scala 64:117 Rename.scala 64:117]
  wire [2:0] _GEN_36 = 5'h4 == io_rob_commit_1_bits_commit_addr ? map_table_4 : _GEN_35; // @[Rename.scala 64:117 Rename.scala 64:117]
  wire [2:0] _GEN_37 = 5'h5 == io_rob_commit_1_bits_commit_addr ? map_table_5 : _GEN_36; // @[Rename.scala 64:117 Rename.scala 64:117]
  wire [2:0] _GEN_38 = 5'h6 == io_rob_commit_1_bits_commit_addr ? map_table_6 : _GEN_37; // @[Rename.scala 64:117 Rename.scala 64:117]
  wire [2:0] _GEN_39 = 5'h7 == io_rob_commit_1_bits_commit_addr ? map_table_7 : _GEN_38; // @[Rename.scala 64:117 Rename.scala 64:117]
  wire [2:0] _GEN_40 = 5'h8 == io_rob_commit_1_bits_commit_addr ? map_table_8 : _GEN_39; // @[Rename.scala 64:117 Rename.scala 64:117]
  wire [2:0] _GEN_41 = 5'h9 == io_rob_commit_1_bits_commit_addr ? map_table_9 : _GEN_40; // @[Rename.scala 64:117 Rename.scala 64:117]
  wire [2:0] _GEN_42 = 5'ha == io_rob_commit_1_bits_commit_addr ? map_table_10 : _GEN_41; // @[Rename.scala 64:117 Rename.scala 64:117]
  wire [2:0] _GEN_43 = 5'hb == io_rob_commit_1_bits_commit_addr ? map_table_11 : _GEN_42; // @[Rename.scala 64:117 Rename.scala 64:117]
  wire [2:0] _GEN_44 = 5'hc == io_rob_commit_1_bits_commit_addr ? map_table_12 : _GEN_43; // @[Rename.scala 64:117 Rename.scala 64:117]
  wire [2:0] _GEN_45 = 5'hd == io_rob_commit_1_bits_commit_addr ? map_table_13 : _GEN_44; // @[Rename.scala 64:117 Rename.scala 64:117]
  wire [2:0] _GEN_46 = 5'he == io_rob_commit_1_bits_commit_addr ? map_table_14 : _GEN_45; // @[Rename.scala 64:117 Rename.scala 64:117]
  wire [2:0] _GEN_47 = 5'hf == io_rob_commit_1_bits_commit_addr ? map_table_15 : _GEN_46; // @[Rename.scala 64:117 Rename.scala 64:117]
  wire [2:0] _GEN_48 = 5'h10 == io_rob_commit_1_bits_commit_addr ? map_table_16 : _GEN_47; // @[Rename.scala 64:117 Rename.scala 64:117]
  wire [2:0] _GEN_49 = 5'h11 == io_rob_commit_1_bits_commit_addr ? map_table_17 : _GEN_48; // @[Rename.scala 64:117 Rename.scala 64:117]
  wire [2:0] _GEN_50 = 5'h12 == io_rob_commit_1_bits_commit_addr ? map_table_18 : _GEN_49; // @[Rename.scala 64:117 Rename.scala 64:117]
  wire [2:0] _GEN_51 = 5'h13 == io_rob_commit_1_bits_commit_addr ? map_table_19 : _GEN_50; // @[Rename.scala 64:117 Rename.scala 64:117]
  wire [2:0] _GEN_52 = 5'h14 == io_rob_commit_1_bits_commit_addr ? map_table_20 : _GEN_51; // @[Rename.scala 64:117 Rename.scala 64:117]
  wire [2:0] _GEN_53 = 5'h15 == io_rob_commit_1_bits_commit_addr ? map_table_21 : _GEN_52; // @[Rename.scala 64:117 Rename.scala 64:117]
  wire [2:0] _GEN_54 = 5'h16 == io_rob_commit_1_bits_commit_addr ? map_table_22 : _GEN_53; // @[Rename.scala 64:117 Rename.scala 64:117]
  wire [2:0] _GEN_55 = 5'h17 == io_rob_commit_1_bits_commit_addr ? map_table_23 : _GEN_54; // @[Rename.scala 64:117 Rename.scala 64:117]
  wire [2:0] _GEN_56 = 5'h18 == io_rob_commit_1_bits_commit_addr ? map_table_24 : _GEN_55; // @[Rename.scala 64:117 Rename.scala 64:117]
  wire [2:0] _GEN_57 = 5'h19 == io_rob_commit_1_bits_commit_addr ? map_table_25 : _GEN_56; // @[Rename.scala 64:117 Rename.scala 64:117]
  wire [2:0] _GEN_58 = 5'h1a == io_rob_commit_1_bits_commit_addr ? map_table_26 : _GEN_57; // @[Rename.scala 64:117 Rename.scala 64:117]
  wire [2:0] _GEN_59 = 5'h1b == io_rob_commit_1_bits_commit_addr ? map_table_27 : _GEN_58; // @[Rename.scala 64:117 Rename.scala 64:117]
  wire [2:0] _GEN_60 = 5'h1c == io_rob_commit_1_bits_commit_addr ? map_table_28 : _GEN_59; // @[Rename.scala 64:117 Rename.scala 64:117]
  wire [2:0] _GEN_61 = 5'h1d == io_rob_commit_1_bits_commit_addr ? map_table_29 : _GEN_60; // @[Rename.scala 64:117 Rename.scala 64:117]
  wire [2:0] _GEN_62 = 5'h1e == io_rob_commit_1_bits_commit_addr ? map_table_30 : _GEN_61; // @[Rename.scala 64:117 Rename.scala 64:117]
  wire [2:0] _GEN_63 = 5'h1f == io_rob_commit_1_bits_commit_addr ? map_table_31 : _GEN_62; // @[Rename.scala 64:117 Rename.scala 64:117]
  wire  _busy_table_wb_T_8 = io_rob_commit_1_valid & io_rob_commit_1_bits_des_rob == _GEN_63; // @[Rename.scala 64:101]
  wire [31:0] _busy_table_wb_T_10 = _busy_table_wb_T_8 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _busy_table_wb_T_11 = _busy_table_wb_T_6 & _busy_table_wb_T_10; // @[Rename.scala 64:85]
  wire [31:0] _busy_table_wb_T_12 = _busy_table_wb_T_5 | _busy_table_wb_T_11; // @[Rename.scala 64:160]
  wire [31:0] _busy_table_wb_T_13 = ~_busy_table_wb_T_12; // @[Rename.scala 64:164]
  wire [31:0] _busy_table_wb_T_14 = busy_table & _busy_table_wb_T_13; // @[Rename.scala 64:34]
  wire [31:0] busy_table_wb = _busy_table_wb_T_14 & 32'hfffffffe; // @[Rename.scala 64:176]
  wire [31:0] busy_table_next = will_busy | busy_table_wb; // @[Rename.scala 65:35]
  reg  rob_init_info_0_is_valid; // @[Rename.scala 73:26]
  reg [2:0] rob_init_info_0_des_rob; // @[Rename.scala 73:26]
  reg [2:0] rob_init_info_0_op1_rob; // @[Rename.scala 73:26]
  reg [2:0] rob_init_info_0_op2_rob; // @[Rename.scala 73:26]
  reg [31:0] rob_init_info_0_op1_regData; // @[Rename.scala 73:26]
  reg [31:0] rob_init_info_0_op2_regData; // @[Rename.scala 73:26]
  reg  rob_init_info_0_op1_in_rob; // @[Rename.scala 73:26]
  reg  rob_init_info_0_op2_in_rob; // @[Rename.scala 73:26]
  reg  rob_init_info_1_is_valid; // @[Rename.scala 73:26]
  reg [2:0] rob_init_info_1_des_rob; // @[Rename.scala 73:26]
  reg [2:0] rob_init_info_1_op1_rob; // @[Rename.scala 73:26]
  reg [2:0] rob_init_info_1_op2_rob; // @[Rename.scala 73:26]
  reg [31:0] rob_init_info_1_op1_regData; // @[Rename.scala 73:26]
  reg [31:0] rob_init_info_1_op2_regData; // @[Rename.scala 73:26]
  reg  rob_init_info_1_op1_in_rob; // @[Rename.scala 73:26]
  reg  rob_init_info_1_op2_in_rob; // @[Rename.scala 73:26]
  reg  rob_init_info_valid; // @[Rename.scala 74:36]
  wire [2:0] _GEN_65 = 5'h1 == io_rename_info_bits_0_op1_addr ? map_table_1 : 3'h0; // @[Rename.scala 79:30 Rename.scala 79:30]
  wire [2:0] _GEN_66 = 5'h2 == io_rename_info_bits_0_op1_addr ? map_table_2 : _GEN_65; // @[Rename.scala 79:30 Rename.scala 79:30]
  wire [2:0] _GEN_67 = 5'h3 == io_rename_info_bits_0_op1_addr ? map_table_3 : _GEN_66; // @[Rename.scala 79:30 Rename.scala 79:30]
  wire [2:0] _GEN_68 = 5'h4 == io_rename_info_bits_0_op1_addr ? map_table_4 : _GEN_67; // @[Rename.scala 79:30 Rename.scala 79:30]
  wire [2:0] _GEN_69 = 5'h5 == io_rename_info_bits_0_op1_addr ? map_table_5 : _GEN_68; // @[Rename.scala 79:30 Rename.scala 79:30]
  wire [2:0] _GEN_70 = 5'h6 == io_rename_info_bits_0_op1_addr ? map_table_6 : _GEN_69; // @[Rename.scala 79:30 Rename.scala 79:30]
  wire [2:0] _GEN_71 = 5'h7 == io_rename_info_bits_0_op1_addr ? map_table_7 : _GEN_70; // @[Rename.scala 79:30 Rename.scala 79:30]
  wire [2:0] _GEN_72 = 5'h8 == io_rename_info_bits_0_op1_addr ? map_table_8 : _GEN_71; // @[Rename.scala 79:30 Rename.scala 79:30]
  wire [2:0] _GEN_73 = 5'h9 == io_rename_info_bits_0_op1_addr ? map_table_9 : _GEN_72; // @[Rename.scala 79:30 Rename.scala 79:30]
  wire [2:0] _GEN_74 = 5'ha == io_rename_info_bits_0_op1_addr ? map_table_10 : _GEN_73; // @[Rename.scala 79:30 Rename.scala 79:30]
  wire [2:0] _GEN_75 = 5'hb == io_rename_info_bits_0_op1_addr ? map_table_11 : _GEN_74; // @[Rename.scala 79:30 Rename.scala 79:30]
  wire [2:0] _GEN_76 = 5'hc == io_rename_info_bits_0_op1_addr ? map_table_12 : _GEN_75; // @[Rename.scala 79:30 Rename.scala 79:30]
  wire [2:0] _GEN_77 = 5'hd == io_rename_info_bits_0_op1_addr ? map_table_13 : _GEN_76; // @[Rename.scala 79:30 Rename.scala 79:30]
  wire [2:0] _GEN_78 = 5'he == io_rename_info_bits_0_op1_addr ? map_table_14 : _GEN_77; // @[Rename.scala 79:30 Rename.scala 79:30]
  wire [2:0] _GEN_79 = 5'hf == io_rename_info_bits_0_op1_addr ? map_table_15 : _GEN_78; // @[Rename.scala 79:30 Rename.scala 79:30]
  wire [2:0] _GEN_80 = 5'h10 == io_rename_info_bits_0_op1_addr ? map_table_16 : _GEN_79; // @[Rename.scala 79:30 Rename.scala 79:30]
  wire [2:0] _GEN_81 = 5'h11 == io_rename_info_bits_0_op1_addr ? map_table_17 : _GEN_80; // @[Rename.scala 79:30 Rename.scala 79:30]
  wire [2:0] _GEN_82 = 5'h12 == io_rename_info_bits_0_op1_addr ? map_table_18 : _GEN_81; // @[Rename.scala 79:30 Rename.scala 79:30]
  wire [2:0] _GEN_83 = 5'h13 == io_rename_info_bits_0_op1_addr ? map_table_19 : _GEN_82; // @[Rename.scala 79:30 Rename.scala 79:30]
  wire [2:0] _GEN_84 = 5'h14 == io_rename_info_bits_0_op1_addr ? map_table_20 : _GEN_83; // @[Rename.scala 79:30 Rename.scala 79:30]
  wire [2:0] _GEN_85 = 5'h15 == io_rename_info_bits_0_op1_addr ? map_table_21 : _GEN_84; // @[Rename.scala 79:30 Rename.scala 79:30]
  wire [2:0] _GEN_86 = 5'h16 == io_rename_info_bits_0_op1_addr ? map_table_22 : _GEN_85; // @[Rename.scala 79:30 Rename.scala 79:30]
  wire [2:0] _GEN_87 = 5'h17 == io_rename_info_bits_0_op1_addr ? map_table_23 : _GEN_86; // @[Rename.scala 79:30 Rename.scala 79:30]
  wire [2:0] _GEN_88 = 5'h18 == io_rename_info_bits_0_op1_addr ? map_table_24 : _GEN_87; // @[Rename.scala 79:30 Rename.scala 79:30]
  wire [2:0] _GEN_89 = 5'h19 == io_rename_info_bits_0_op1_addr ? map_table_25 : _GEN_88; // @[Rename.scala 79:30 Rename.scala 79:30]
  wire [2:0] _GEN_90 = 5'h1a == io_rename_info_bits_0_op1_addr ? map_table_26 : _GEN_89; // @[Rename.scala 79:30 Rename.scala 79:30]
  wire [2:0] _GEN_91 = 5'h1b == io_rename_info_bits_0_op1_addr ? map_table_27 : _GEN_90; // @[Rename.scala 79:30 Rename.scala 79:30]
  wire [2:0] _GEN_92 = 5'h1c == io_rename_info_bits_0_op1_addr ? map_table_28 : _GEN_91; // @[Rename.scala 79:30 Rename.scala 79:30]
  wire [2:0] _GEN_93 = 5'h1d == io_rename_info_bits_0_op1_addr ? map_table_29 : _GEN_92; // @[Rename.scala 79:30 Rename.scala 79:30]
  wire [2:0] _GEN_97 = 5'h1 == io_rename_info_bits_0_op2_addr ? map_table_1 : 3'h0; // @[Rename.scala 82:30 Rename.scala 82:30]
  wire [2:0] _GEN_98 = 5'h2 == io_rename_info_bits_0_op2_addr ? map_table_2 : _GEN_97; // @[Rename.scala 82:30 Rename.scala 82:30]
  wire [2:0] _GEN_99 = 5'h3 == io_rename_info_bits_0_op2_addr ? map_table_3 : _GEN_98; // @[Rename.scala 82:30 Rename.scala 82:30]
  wire [2:0] _GEN_100 = 5'h4 == io_rename_info_bits_0_op2_addr ? map_table_4 : _GEN_99; // @[Rename.scala 82:30 Rename.scala 82:30]
  wire [2:0] _GEN_101 = 5'h5 == io_rename_info_bits_0_op2_addr ? map_table_5 : _GEN_100; // @[Rename.scala 82:30 Rename.scala 82:30]
  wire [2:0] _GEN_102 = 5'h6 == io_rename_info_bits_0_op2_addr ? map_table_6 : _GEN_101; // @[Rename.scala 82:30 Rename.scala 82:30]
  wire [2:0] _GEN_103 = 5'h7 == io_rename_info_bits_0_op2_addr ? map_table_7 : _GEN_102; // @[Rename.scala 82:30 Rename.scala 82:30]
  wire [2:0] _GEN_104 = 5'h8 == io_rename_info_bits_0_op2_addr ? map_table_8 : _GEN_103; // @[Rename.scala 82:30 Rename.scala 82:30]
  wire [2:0] _GEN_105 = 5'h9 == io_rename_info_bits_0_op2_addr ? map_table_9 : _GEN_104; // @[Rename.scala 82:30 Rename.scala 82:30]
  wire [2:0] _GEN_106 = 5'ha == io_rename_info_bits_0_op2_addr ? map_table_10 : _GEN_105; // @[Rename.scala 82:30 Rename.scala 82:30]
  wire [2:0] _GEN_107 = 5'hb == io_rename_info_bits_0_op2_addr ? map_table_11 : _GEN_106; // @[Rename.scala 82:30 Rename.scala 82:30]
  wire [2:0] _GEN_108 = 5'hc == io_rename_info_bits_0_op2_addr ? map_table_12 : _GEN_107; // @[Rename.scala 82:30 Rename.scala 82:30]
  wire [2:0] _GEN_109 = 5'hd == io_rename_info_bits_0_op2_addr ? map_table_13 : _GEN_108; // @[Rename.scala 82:30 Rename.scala 82:30]
  wire [2:0] _GEN_110 = 5'he == io_rename_info_bits_0_op2_addr ? map_table_14 : _GEN_109; // @[Rename.scala 82:30 Rename.scala 82:30]
  wire [2:0] _GEN_111 = 5'hf == io_rename_info_bits_0_op2_addr ? map_table_15 : _GEN_110; // @[Rename.scala 82:30 Rename.scala 82:30]
  wire [2:0] _GEN_112 = 5'h10 == io_rename_info_bits_0_op2_addr ? map_table_16 : _GEN_111; // @[Rename.scala 82:30 Rename.scala 82:30]
  wire [2:0] _GEN_113 = 5'h11 == io_rename_info_bits_0_op2_addr ? map_table_17 : _GEN_112; // @[Rename.scala 82:30 Rename.scala 82:30]
  wire [2:0] _GEN_114 = 5'h12 == io_rename_info_bits_0_op2_addr ? map_table_18 : _GEN_113; // @[Rename.scala 82:30 Rename.scala 82:30]
  wire [2:0] _GEN_115 = 5'h13 == io_rename_info_bits_0_op2_addr ? map_table_19 : _GEN_114; // @[Rename.scala 82:30 Rename.scala 82:30]
  wire [2:0] _GEN_116 = 5'h14 == io_rename_info_bits_0_op2_addr ? map_table_20 : _GEN_115; // @[Rename.scala 82:30 Rename.scala 82:30]
  wire [2:0] _GEN_117 = 5'h15 == io_rename_info_bits_0_op2_addr ? map_table_21 : _GEN_116; // @[Rename.scala 82:30 Rename.scala 82:30]
  wire [2:0] _GEN_118 = 5'h16 == io_rename_info_bits_0_op2_addr ? map_table_22 : _GEN_117; // @[Rename.scala 82:30 Rename.scala 82:30]
  wire [2:0] _GEN_119 = 5'h17 == io_rename_info_bits_0_op2_addr ? map_table_23 : _GEN_118; // @[Rename.scala 82:30 Rename.scala 82:30]
  wire [2:0] _GEN_120 = 5'h18 == io_rename_info_bits_0_op2_addr ? map_table_24 : _GEN_119; // @[Rename.scala 82:30 Rename.scala 82:30]
  wire [2:0] _GEN_121 = 5'h19 == io_rename_info_bits_0_op2_addr ? map_table_25 : _GEN_120; // @[Rename.scala 82:30 Rename.scala 82:30]
  wire [2:0] _GEN_122 = 5'h1a == io_rename_info_bits_0_op2_addr ? map_table_26 : _GEN_121; // @[Rename.scala 82:30 Rename.scala 82:30]
  wire [2:0] _GEN_123 = 5'h1b == io_rename_info_bits_0_op2_addr ? map_table_27 : _GEN_122; // @[Rename.scala 82:30 Rename.scala 82:30]
  wire [2:0] _GEN_124 = 5'h1c == io_rename_info_bits_0_op2_addr ? map_table_28 : _GEN_123; // @[Rename.scala 82:30 Rename.scala 82:30]
  wire [2:0] _GEN_125 = 5'h1d == io_rename_info_bits_0_op2_addr ? map_table_29 : _GEN_124; // @[Rename.scala 82:30 Rename.scala 82:30]
  wire [31:0] _rob_init_info_0_op1_in_rob_T = busy_table_wb >> io_rename_info_bits_0_op1_addr; // @[Rename.scala 85:221]
  wire [31:0] _rob_init_info_0_op2_in_rob_T = busy_table_wb >> io_rename_info_bits_0_op2_addr; // @[Rename.scala 86:221]
  wire  _rob_init_info_1_op1_rob_T_1 = io_rename_info_bits_0_is_valid & io_rename_info_bits_0_des_addr ==
    io_rename_info_bits_1_op1_addr; // @[Rename.scala 80:53]
  wire [2:0] _GEN_129 = 5'h1 == io_rename_info_bits_1_op1_addr ? map_table_1 : 3'h0; // @[Rename.scala 80:20 Rename.scala 80:20]
  wire [2:0] _GEN_130 = 5'h2 == io_rename_info_bits_1_op1_addr ? map_table_2 : _GEN_129; // @[Rename.scala 80:20 Rename.scala 80:20]
  wire [2:0] _GEN_131 = 5'h3 == io_rename_info_bits_1_op1_addr ? map_table_3 : _GEN_130; // @[Rename.scala 80:20 Rename.scala 80:20]
  wire [2:0] _GEN_132 = 5'h4 == io_rename_info_bits_1_op1_addr ? map_table_4 : _GEN_131; // @[Rename.scala 80:20 Rename.scala 80:20]
  wire [2:0] _GEN_133 = 5'h5 == io_rename_info_bits_1_op1_addr ? map_table_5 : _GEN_132; // @[Rename.scala 80:20 Rename.scala 80:20]
  wire [2:0] _GEN_134 = 5'h6 == io_rename_info_bits_1_op1_addr ? map_table_6 : _GEN_133; // @[Rename.scala 80:20 Rename.scala 80:20]
  wire [2:0] _GEN_135 = 5'h7 == io_rename_info_bits_1_op1_addr ? map_table_7 : _GEN_134; // @[Rename.scala 80:20 Rename.scala 80:20]
  wire [2:0] _GEN_136 = 5'h8 == io_rename_info_bits_1_op1_addr ? map_table_8 : _GEN_135; // @[Rename.scala 80:20 Rename.scala 80:20]
  wire [2:0] _GEN_137 = 5'h9 == io_rename_info_bits_1_op1_addr ? map_table_9 : _GEN_136; // @[Rename.scala 80:20 Rename.scala 80:20]
  wire [2:0] _GEN_138 = 5'ha == io_rename_info_bits_1_op1_addr ? map_table_10 : _GEN_137; // @[Rename.scala 80:20 Rename.scala 80:20]
  wire [2:0] _GEN_139 = 5'hb == io_rename_info_bits_1_op1_addr ? map_table_11 : _GEN_138; // @[Rename.scala 80:20 Rename.scala 80:20]
  wire [2:0] _GEN_140 = 5'hc == io_rename_info_bits_1_op1_addr ? map_table_12 : _GEN_139; // @[Rename.scala 80:20 Rename.scala 80:20]
  wire [2:0] _GEN_141 = 5'hd == io_rename_info_bits_1_op1_addr ? map_table_13 : _GEN_140; // @[Rename.scala 80:20 Rename.scala 80:20]
  wire [2:0] _GEN_142 = 5'he == io_rename_info_bits_1_op1_addr ? map_table_14 : _GEN_141; // @[Rename.scala 80:20 Rename.scala 80:20]
  wire [2:0] _GEN_143 = 5'hf == io_rename_info_bits_1_op1_addr ? map_table_15 : _GEN_142; // @[Rename.scala 80:20 Rename.scala 80:20]
  wire [2:0] _GEN_144 = 5'h10 == io_rename_info_bits_1_op1_addr ? map_table_16 : _GEN_143; // @[Rename.scala 80:20 Rename.scala 80:20]
  wire [2:0] _GEN_145 = 5'h11 == io_rename_info_bits_1_op1_addr ? map_table_17 : _GEN_144; // @[Rename.scala 80:20 Rename.scala 80:20]
  wire [2:0] _GEN_146 = 5'h12 == io_rename_info_bits_1_op1_addr ? map_table_18 : _GEN_145; // @[Rename.scala 80:20 Rename.scala 80:20]
  wire [2:0] _GEN_147 = 5'h13 == io_rename_info_bits_1_op1_addr ? map_table_19 : _GEN_146; // @[Rename.scala 80:20 Rename.scala 80:20]
  wire [2:0] _GEN_148 = 5'h14 == io_rename_info_bits_1_op1_addr ? map_table_20 : _GEN_147; // @[Rename.scala 80:20 Rename.scala 80:20]
  wire [2:0] _GEN_149 = 5'h15 == io_rename_info_bits_1_op1_addr ? map_table_21 : _GEN_148; // @[Rename.scala 80:20 Rename.scala 80:20]
  wire [2:0] _GEN_150 = 5'h16 == io_rename_info_bits_1_op1_addr ? map_table_22 : _GEN_149; // @[Rename.scala 80:20 Rename.scala 80:20]
  wire [2:0] _GEN_151 = 5'h17 == io_rename_info_bits_1_op1_addr ? map_table_23 : _GEN_150; // @[Rename.scala 80:20 Rename.scala 80:20]
  wire [2:0] _GEN_152 = 5'h18 == io_rename_info_bits_1_op1_addr ? map_table_24 : _GEN_151; // @[Rename.scala 80:20 Rename.scala 80:20]
  wire [2:0] _GEN_153 = 5'h19 == io_rename_info_bits_1_op1_addr ? map_table_25 : _GEN_152; // @[Rename.scala 80:20 Rename.scala 80:20]
  wire [2:0] _GEN_154 = 5'h1a == io_rename_info_bits_1_op1_addr ? map_table_26 : _GEN_153; // @[Rename.scala 80:20 Rename.scala 80:20]
  wire [2:0] _GEN_155 = 5'h1b == io_rename_info_bits_1_op1_addr ? map_table_27 : _GEN_154; // @[Rename.scala 80:20 Rename.scala 80:20]
  wire [2:0] _GEN_156 = 5'h1c == io_rename_info_bits_1_op1_addr ? map_table_28 : _GEN_155; // @[Rename.scala 80:20 Rename.scala 80:20]
  wire [2:0] _GEN_157 = 5'h1d == io_rename_info_bits_1_op1_addr ? map_table_29 : _GEN_156; // @[Rename.scala 80:20 Rename.scala 80:20]
  wire [2:0] _GEN_158 = 5'h1e == io_rename_info_bits_1_op1_addr ? map_table_30 : _GEN_157; // @[Rename.scala 80:20 Rename.scala 80:20]
  wire  _rob_init_info_1_op2_rob_T_1 = io_rename_info_bits_0_is_valid & io_rename_info_bits_0_des_addr ==
    io_rename_info_bits_1_op2_addr; // @[Rename.scala 83:53]
  wire [2:0] _GEN_161 = 5'h1 == io_rename_info_bits_1_op2_addr ? map_table_1 : 3'h0; // @[Rename.scala 83:20 Rename.scala 83:20]
  wire [2:0] _GEN_162 = 5'h2 == io_rename_info_bits_1_op2_addr ? map_table_2 : _GEN_161; // @[Rename.scala 83:20 Rename.scala 83:20]
  wire [2:0] _GEN_163 = 5'h3 == io_rename_info_bits_1_op2_addr ? map_table_3 : _GEN_162; // @[Rename.scala 83:20 Rename.scala 83:20]
  wire [2:0] _GEN_164 = 5'h4 == io_rename_info_bits_1_op2_addr ? map_table_4 : _GEN_163; // @[Rename.scala 83:20 Rename.scala 83:20]
  wire [2:0] _GEN_165 = 5'h5 == io_rename_info_bits_1_op2_addr ? map_table_5 : _GEN_164; // @[Rename.scala 83:20 Rename.scala 83:20]
  wire [2:0] _GEN_166 = 5'h6 == io_rename_info_bits_1_op2_addr ? map_table_6 : _GEN_165; // @[Rename.scala 83:20 Rename.scala 83:20]
  wire [2:0] _GEN_167 = 5'h7 == io_rename_info_bits_1_op2_addr ? map_table_7 : _GEN_166; // @[Rename.scala 83:20 Rename.scala 83:20]
  wire [2:0] _GEN_168 = 5'h8 == io_rename_info_bits_1_op2_addr ? map_table_8 : _GEN_167; // @[Rename.scala 83:20 Rename.scala 83:20]
  wire [2:0] _GEN_169 = 5'h9 == io_rename_info_bits_1_op2_addr ? map_table_9 : _GEN_168; // @[Rename.scala 83:20 Rename.scala 83:20]
  wire [2:0] _GEN_170 = 5'ha == io_rename_info_bits_1_op2_addr ? map_table_10 : _GEN_169; // @[Rename.scala 83:20 Rename.scala 83:20]
  wire [2:0] _GEN_171 = 5'hb == io_rename_info_bits_1_op2_addr ? map_table_11 : _GEN_170; // @[Rename.scala 83:20 Rename.scala 83:20]
  wire [2:0] _GEN_172 = 5'hc == io_rename_info_bits_1_op2_addr ? map_table_12 : _GEN_171; // @[Rename.scala 83:20 Rename.scala 83:20]
  wire [2:0] _GEN_173 = 5'hd == io_rename_info_bits_1_op2_addr ? map_table_13 : _GEN_172; // @[Rename.scala 83:20 Rename.scala 83:20]
  wire [2:0] _GEN_174 = 5'he == io_rename_info_bits_1_op2_addr ? map_table_14 : _GEN_173; // @[Rename.scala 83:20 Rename.scala 83:20]
  wire [2:0] _GEN_175 = 5'hf == io_rename_info_bits_1_op2_addr ? map_table_15 : _GEN_174; // @[Rename.scala 83:20 Rename.scala 83:20]
  wire [2:0] _GEN_176 = 5'h10 == io_rename_info_bits_1_op2_addr ? map_table_16 : _GEN_175; // @[Rename.scala 83:20 Rename.scala 83:20]
  wire [2:0] _GEN_177 = 5'h11 == io_rename_info_bits_1_op2_addr ? map_table_17 : _GEN_176; // @[Rename.scala 83:20 Rename.scala 83:20]
  wire [2:0] _GEN_178 = 5'h12 == io_rename_info_bits_1_op2_addr ? map_table_18 : _GEN_177; // @[Rename.scala 83:20 Rename.scala 83:20]
  wire [2:0] _GEN_179 = 5'h13 == io_rename_info_bits_1_op2_addr ? map_table_19 : _GEN_178; // @[Rename.scala 83:20 Rename.scala 83:20]
  wire [2:0] _GEN_180 = 5'h14 == io_rename_info_bits_1_op2_addr ? map_table_20 : _GEN_179; // @[Rename.scala 83:20 Rename.scala 83:20]
  wire [2:0] _GEN_181 = 5'h15 == io_rename_info_bits_1_op2_addr ? map_table_21 : _GEN_180; // @[Rename.scala 83:20 Rename.scala 83:20]
  wire [2:0] _GEN_182 = 5'h16 == io_rename_info_bits_1_op2_addr ? map_table_22 : _GEN_181; // @[Rename.scala 83:20 Rename.scala 83:20]
  wire [2:0] _GEN_183 = 5'h17 == io_rename_info_bits_1_op2_addr ? map_table_23 : _GEN_182; // @[Rename.scala 83:20 Rename.scala 83:20]
  wire [2:0] _GEN_184 = 5'h18 == io_rename_info_bits_1_op2_addr ? map_table_24 : _GEN_183; // @[Rename.scala 83:20 Rename.scala 83:20]
  wire [2:0] _GEN_185 = 5'h19 == io_rename_info_bits_1_op2_addr ? map_table_25 : _GEN_184; // @[Rename.scala 83:20 Rename.scala 83:20]
  wire [2:0] _GEN_186 = 5'h1a == io_rename_info_bits_1_op2_addr ? map_table_26 : _GEN_185; // @[Rename.scala 83:20 Rename.scala 83:20]
  wire [2:0] _GEN_187 = 5'h1b == io_rename_info_bits_1_op2_addr ? map_table_27 : _GEN_186; // @[Rename.scala 83:20 Rename.scala 83:20]
  wire [2:0] _GEN_188 = 5'h1c == io_rename_info_bits_1_op2_addr ? map_table_28 : _GEN_187; // @[Rename.scala 83:20 Rename.scala 83:20]
  wire [2:0] _GEN_189 = 5'h1d == io_rename_info_bits_1_op2_addr ? map_table_29 : _GEN_188; // @[Rename.scala 83:20 Rename.scala 83:20]
  wire [2:0] _GEN_190 = 5'h1e == io_rename_info_bits_1_op2_addr ? map_table_30 : _GEN_189; // @[Rename.scala 83:20 Rename.scala 83:20]
  wire  _rob_init_info_1_op1_in_rob_T_2 = io_rename_info_bits_0_des_addr != 5'h0; // @[Rename.scala 85:190]
  wire [31:0] _rob_init_info_1_op1_in_rob_T_4 = busy_table_wb >> io_rename_info_bits_1_op1_addr; // @[Rename.scala 85:221]
  wire [31:0] _rob_init_info_1_op2_in_rob_T_4 = busy_table_wb >> io_rename_info_bits_1_op2_addr; // @[Rename.scala 86:221]
  assign io_reg_read_0_op1_addr = io_rename_info_bits_0_op1_addr; // @[Rename.scala 87:29]
  assign io_reg_read_0_op2_addr = io_rename_info_bits_0_op2_addr; // @[Rename.scala 88:29]
  assign io_reg_read_1_op1_addr = io_rename_info_bits_1_op1_addr; // @[Rename.scala 87:29]
  assign io_reg_read_1_op2_addr = io_rename_info_bits_1_op2_addr; // @[Rename.scala 88:29]
  assign io_rob_init_info_valid = rob_init_info_valid; // @[Rename.scala 76:26]
  assign io_rob_init_info_bits_0_is_valid = rob_init_info_0_is_valid; // @[Rename.scala 75:25]
  assign io_rob_init_info_bits_0_des_rob = rob_init_info_0_des_rob; // @[Rename.scala 75:25]
  assign io_rob_init_info_bits_0_op1_rob = rob_init_info_0_op1_rob; // @[Rename.scala 75:25]
  assign io_rob_init_info_bits_0_op2_rob = rob_init_info_0_op2_rob; // @[Rename.scala 75:25]
  assign io_rob_init_info_bits_0_op1_regData = rob_init_info_0_op1_regData; // @[Rename.scala 75:25]
  assign io_rob_init_info_bits_0_op2_regData = rob_init_info_0_op2_regData; // @[Rename.scala 75:25]
  assign io_rob_init_info_bits_0_op1_in_rob = rob_init_info_0_op1_in_rob; // @[Rename.scala 75:25]
  assign io_rob_init_info_bits_0_op2_in_rob = rob_init_info_0_op2_in_rob; // @[Rename.scala 75:25]
  assign io_rob_init_info_bits_1_is_valid = rob_init_info_1_is_valid; // @[Rename.scala 75:25]
  assign io_rob_init_info_bits_1_des_rob = rob_init_info_1_des_rob; // @[Rename.scala 75:25]
  assign io_rob_init_info_bits_1_op1_rob = rob_init_info_1_op1_rob; // @[Rename.scala 75:25]
  assign io_rob_init_info_bits_1_op2_rob = rob_init_info_1_op2_rob; // @[Rename.scala 75:25]
  assign io_rob_init_info_bits_1_op1_regData = rob_init_info_1_op1_regData; // @[Rename.scala 75:25]
  assign io_rob_init_info_bits_1_op2_regData = rob_init_info_1_op2_regData; // @[Rename.scala 75:25]
  assign io_rob_init_info_bits_1_op1_in_rob = rob_init_info_1_op1_in_rob; // @[Rename.scala 75:25]
  assign io_rob_init_info_bits_1_op2_in_rob = rob_init_info_1_op2_in_rob; // @[Rename.scala 75:25]
  always @(posedge clock) begin
    if (reset) begin // @[Rename.scala 60:27]
      busy_table <= 32'h0; // @[Rename.scala 60:27]
    end else if (io_need_flush) begin // @[Rename.scala 66:18]
      busy_table <= 32'h0;
    end else begin
      busy_table <= busy_table_next;
    end
    if (reset) begin // @[Rename.scala 61:26]
      map_table_1 <= 3'h0; // @[Rename.scala 61:26]
    end else if (_will_busy_T_6 & _will_busy_T_5[1]) begin // @[Rename.scala 70:101]
      map_table_1 <= io_rename_info_bits_1_des_rob;
    end else if (_will_busy_T_1 & _will_busy_T[1]) begin // @[Rename.scala 70:101]
      map_table_1 <= io_rename_info_bits_0_des_rob;
    end
    if (reset) begin // @[Rename.scala 61:26]
      map_table_2 <= 3'h0; // @[Rename.scala 61:26]
    end else if (_will_busy_T_6 & _will_busy_T_5[2]) begin // @[Rename.scala 70:101]
      map_table_2 <= io_rename_info_bits_1_des_rob;
    end else if (_will_busy_T_1 & _will_busy_T[2]) begin // @[Rename.scala 70:101]
      map_table_2 <= io_rename_info_bits_0_des_rob;
    end
    if (reset) begin // @[Rename.scala 61:26]
      map_table_3 <= 3'h0; // @[Rename.scala 61:26]
    end else if (_will_busy_T_6 & _will_busy_T_5[3]) begin // @[Rename.scala 70:101]
      map_table_3 <= io_rename_info_bits_1_des_rob;
    end else if (_will_busy_T_1 & _will_busy_T[3]) begin // @[Rename.scala 70:101]
      map_table_3 <= io_rename_info_bits_0_des_rob;
    end
    if (reset) begin // @[Rename.scala 61:26]
      map_table_4 <= 3'h0; // @[Rename.scala 61:26]
    end else if (_will_busy_T_6 & _will_busy_T_5[4]) begin // @[Rename.scala 70:101]
      map_table_4 <= io_rename_info_bits_1_des_rob;
    end else if (_will_busy_T_1 & _will_busy_T[4]) begin // @[Rename.scala 70:101]
      map_table_4 <= io_rename_info_bits_0_des_rob;
    end
    if (reset) begin // @[Rename.scala 61:26]
      map_table_5 <= 3'h0; // @[Rename.scala 61:26]
    end else if (_will_busy_T_6 & _will_busy_T_5[5]) begin // @[Rename.scala 70:101]
      map_table_5 <= io_rename_info_bits_1_des_rob;
    end else if (_will_busy_T_1 & _will_busy_T[5]) begin // @[Rename.scala 70:101]
      map_table_5 <= io_rename_info_bits_0_des_rob;
    end
    if (reset) begin // @[Rename.scala 61:26]
      map_table_6 <= 3'h0; // @[Rename.scala 61:26]
    end else if (_will_busy_T_6 & _will_busy_T_5[6]) begin // @[Rename.scala 70:101]
      map_table_6 <= io_rename_info_bits_1_des_rob;
    end else if (_will_busy_T_1 & _will_busy_T[6]) begin // @[Rename.scala 70:101]
      map_table_6 <= io_rename_info_bits_0_des_rob;
    end
    if (reset) begin // @[Rename.scala 61:26]
      map_table_7 <= 3'h0; // @[Rename.scala 61:26]
    end else if (_will_busy_T_6 & _will_busy_T_5[7]) begin // @[Rename.scala 70:101]
      map_table_7 <= io_rename_info_bits_1_des_rob;
    end else if (_will_busy_T_1 & _will_busy_T[7]) begin // @[Rename.scala 70:101]
      map_table_7 <= io_rename_info_bits_0_des_rob;
    end
    if (reset) begin // @[Rename.scala 61:26]
      map_table_8 <= 3'h0; // @[Rename.scala 61:26]
    end else if (_will_busy_T_6 & _will_busy_T_5[8]) begin // @[Rename.scala 70:101]
      map_table_8 <= io_rename_info_bits_1_des_rob;
    end else if (_will_busy_T_1 & _will_busy_T[8]) begin // @[Rename.scala 70:101]
      map_table_8 <= io_rename_info_bits_0_des_rob;
    end
    if (reset) begin // @[Rename.scala 61:26]
      map_table_9 <= 3'h0; // @[Rename.scala 61:26]
    end else if (_will_busy_T_6 & _will_busy_T_5[9]) begin // @[Rename.scala 70:101]
      map_table_9 <= io_rename_info_bits_1_des_rob;
    end else if (_will_busy_T_1 & _will_busy_T[9]) begin // @[Rename.scala 70:101]
      map_table_9 <= io_rename_info_bits_0_des_rob;
    end
    if (reset) begin // @[Rename.scala 61:26]
      map_table_10 <= 3'h0; // @[Rename.scala 61:26]
    end else if (_will_busy_T_6 & _will_busy_T_5[10]) begin // @[Rename.scala 70:101]
      map_table_10 <= io_rename_info_bits_1_des_rob;
    end else if (_will_busy_T_1 & _will_busy_T[10]) begin // @[Rename.scala 70:101]
      map_table_10 <= io_rename_info_bits_0_des_rob;
    end
    if (reset) begin // @[Rename.scala 61:26]
      map_table_11 <= 3'h0; // @[Rename.scala 61:26]
    end else if (_will_busy_T_6 & _will_busy_T_5[11]) begin // @[Rename.scala 70:101]
      map_table_11 <= io_rename_info_bits_1_des_rob;
    end else if (_will_busy_T_1 & _will_busy_T[11]) begin // @[Rename.scala 70:101]
      map_table_11 <= io_rename_info_bits_0_des_rob;
    end
    if (reset) begin // @[Rename.scala 61:26]
      map_table_12 <= 3'h0; // @[Rename.scala 61:26]
    end else if (_will_busy_T_6 & _will_busy_T_5[12]) begin // @[Rename.scala 70:101]
      map_table_12 <= io_rename_info_bits_1_des_rob;
    end else if (_will_busy_T_1 & _will_busy_T[12]) begin // @[Rename.scala 70:101]
      map_table_12 <= io_rename_info_bits_0_des_rob;
    end
    if (reset) begin // @[Rename.scala 61:26]
      map_table_13 <= 3'h0; // @[Rename.scala 61:26]
    end else if (_will_busy_T_6 & _will_busy_T_5[13]) begin // @[Rename.scala 70:101]
      map_table_13 <= io_rename_info_bits_1_des_rob;
    end else if (_will_busy_T_1 & _will_busy_T[13]) begin // @[Rename.scala 70:101]
      map_table_13 <= io_rename_info_bits_0_des_rob;
    end
    if (reset) begin // @[Rename.scala 61:26]
      map_table_14 <= 3'h0; // @[Rename.scala 61:26]
    end else if (_will_busy_T_6 & _will_busy_T_5[14]) begin // @[Rename.scala 70:101]
      map_table_14 <= io_rename_info_bits_1_des_rob;
    end else if (_will_busy_T_1 & _will_busy_T[14]) begin // @[Rename.scala 70:101]
      map_table_14 <= io_rename_info_bits_0_des_rob;
    end
    if (reset) begin // @[Rename.scala 61:26]
      map_table_15 <= 3'h0; // @[Rename.scala 61:26]
    end else if (_will_busy_T_6 & _will_busy_T_5[15]) begin // @[Rename.scala 70:101]
      map_table_15 <= io_rename_info_bits_1_des_rob;
    end else if (_will_busy_T_1 & _will_busy_T[15]) begin // @[Rename.scala 70:101]
      map_table_15 <= io_rename_info_bits_0_des_rob;
    end
    if (reset) begin // @[Rename.scala 61:26]
      map_table_16 <= 3'h0; // @[Rename.scala 61:26]
    end else if (_will_busy_T_6 & _will_busy_T_5[16]) begin // @[Rename.scala 70:101]
      map_table_16 <= io_rename_info_bits_1_des_rob;
    end else if (_will_busy_T_1 & _will_busy_T[16]) begin // @[Rename.scala 70:101]
      map_table_16 <= io_rename_info_bits_0_des_rob;
    end
    if (reset) begin // @[Rename.scala 61:26]
      map_table_17 <= 3'h0; // @[Rename.scala 61:26]
    end else if (_will_busy_T_6 & _will_busy_T_5[17]) begin // @[Rename.scala 70:101]
      map_table_17 <= io_rename_info_bits_1_des_rob;
    end else if (_will_busy_T_1 & _will_busy_T[17]) begin // @[Rename.scala 70:101]
      map_table_17 <= io_rename_info_bits_0_des_rob;
    end
    if (reset) begin // @[Rename.scala 61:26]
      map_table_18 <= 3'h0; // @[Rename.scala 61:26]
    end else if (_will_busy_T_6 & _will_busy_T_5[18]) begin // @[Rename.scala 70:101]
      map_table_18 <= io_rename_info_bits_1_des_rob;
    end else if (_will_busy_T_1 & _will_busy_T[18]) begin // @[Rename.scala 70:101]
      map_table_18 <= io_rename_info_bits_0_des_rob;
    end
    if (reset) begin // @[Rename.scala 61:26]
      map_table_19 <= 3'h0; // @[Rename.scala 61:26]
    end else if (_will_busy_T_6 & _will_busy_T_5[19]) begin // @[Rename.scala 70:101]
      map_table_19 <= io_rename_info_bits_1_des_rob;
    end else if (_will_busy_T_1 & _will_busy_T[19]) begin // @[Rename.scala 70:101]
      map_table_19 <= io_rename_info_bits_0_des_rob;
    end
    if (reset) begin // @[Rename.scala 61:26]
      map_table_20 <= 3'h0; // @[Rename.scala 61:26]
    end else if (_will_busy_T_6 & _will_busy_T_5[20]) begin // @[Rename.scala 70:101]
      map_table_20 <= io_rename_info_bits_1_des_rob;
    end else if (_will_busy_T_1 & _will_busy_T[20]) begin // @[Rename.scala 70:101]
      map_table_20 <= io_rename_info_bits_0_des_rob;
    end
    if (reset) begin // @[Rename.scala 61:26]
      map_table_21 <= 3'h0; // @[Rename.scala 61:26]
    end else if (_will_busy_T_6 & _will_busy_T_5[21]) begin // @[Rename.scala 70:101]
      map_table_21 <= io_rename_info_bits_1_des_rob;
    end else if (_will_busy_T_1 & _will_busy_T[21]) begin // @[Rename.scala 70:101]
      map_table_21 <= io_rename_info_bits_0_des_rob;
    end
    if (reset) begin // @[Rename.scala 61:26]
      map_table_22 <= 3'h0; // @[Rename.scala 61:26]
    end else if (_will_busy_T_6 & _will_busy_T_5[22]) begin // @[Rename.scala 70:101]
      map_table_22 <= io_rename_info_bits_1_des_rob;
    end else if (_will_busy_T_1 & _will_busy_T[22]) begin // @[Rename.scala 70:101]
      map_table_22 <= io_rename_info_bits_0_des_rob;
    end
    if (reset) begin // @[Rename.scala 61:26]
      map_table_23 <= 3'h0; // @[Rename.scala 61:26]
    end else if (_will_busy_T_6 & _will_busy_T_5[23]) begin // @[Rename.scala 70:101]
      map_table_23 <= io_rename_info_bits_1_des_rob;
    end else if (_will_busy_T_1 & _will_busy_T[23]) begin // @[Rename.scala 70:101]
      map_table_23 <= io_rename_info_bits_0_des_rob;
    end
    if (reset) begin // @[Rename.scala 61:26]
      map_table_24 <= 3'h0; // @[Rename.scala 61:26]
    end else if (_will_busy_T_6 & _will_busy_T_5[24]) begin // @[Rename.scala 70:101]
      map_table_24 <= io_rename_info_bits_1_des_rob;
    end else if (_will_busy_T_1 & _will_busy_T[24]) begin // @[Rename.scala 70:101]
      map_table_24 <= io_rename_info_bits_0_des_rob;
    end
    if (reset) begin // @[Rename.scala 61:26]
      map_table_25 <= 3'h0; // @[Rename.scala 61:26]
    end else if (_will_busy_T_6 & _will_busy_T_5[25]) begin // @[Rename.scala 70:101]
      map_table_25 <= io_rename_info_bits_1_des_rob;
    end else if (_will_busy_T_1 & _will_busy_T[25]) begin // @[Rename.scala 70:101]
      map_table_25 <= io_rename_info_bits_0_des_rob;
    end
    if (reset) begin // @[Rename.scala 61:26]
      map_table_26 <= 3'h0; // @[Rename.scala 61:26]
    end else if (_will_busy_T_6 & _will_busy_T_5[26]) begin // @[Rename.scala 70:101]
      map_table_26 <= io_rename_info_bits_1_des_rob;
    end else if (_will_busy_T_1 & _will_busy_T[26]) begin // @[Rename.scala 70:101]
      map_table_26 <= io_rename_info_bits_0_des_rob;
    end
    if (reset) begin // @[Rename.scala 61:26]
      map_table_27 <= 3'h0; // @[Rename.scala 61:26]
    end else if (_will_busy_T_6 & _will_busy_T_5[27]) begin // @[Rename.scala 70:101]
      map_table_27 <= io_rename_info_bits_1_des_rob;
    end else if (_will_busy_T_1 & _will_busy_T[27]) begin // @[Rename.scala 70:101]
      map_table_27 <= io_rename_info_bits_0_des_rob;
    end
    if (reset) begin // @[Rename.scala 61:26]
      map_table_28 <= 3'h0; // @[Rename.scala 61:26]
    end else if (_will_busy_T_6 & _will_busy_T_5[28]) begin // @[Rename.scala 70:101]
      map_table_28 <= io_rename_info_bits_1_des_rob;
    end else if (_will_busy_T_1 & _will_busy_T[28]) begin // @[Rename.scala 70:101]
      map_table_28 <= io_rename_info_bits_0_des_rob;
    end
    if (reset) begin // @[Rename.scala 61:26]
      map_table_29 <= 3'h0; // @[Rename.scala 61:26]
    end else if (_will_busy_T_6 & _will_busy_T_5[29]) begin // @[Rename.scala 70:101]
      map_table_29 <= io_rename_info_bits_1_des_rob;
    end else if (_will_busy_T_1 & _will_busy_T[29]) begin // @[Rename.scala 70:101]
      map_table_29 <= io_rename_info_bits_0_des_rob;
    end
    if (reset) begin // @[Rename.scala 61:26]
      map_table_30 <= 3'h0; // @[Rename.scala 61:26]
    end else if (_will_busy_T_6 & _will_busy_T_5[30]) begin // @[Rename.scala 70:101]
      map_table_30 <= io_rename_info_bits_1_des_rob;
    end else if (_will_busy_T_1 & _will_busy_T[30]) begin // @[Rename.scala 70:101]
      map_table_30 <= io_rename_info_bits_0_des_rob;
    end
    if (reset) begin // @[Rename.scala 61:26]
      map_table_31 <= 3'h0; // @[Rename.scala 61:26]
    end else if (_will_busy_T_6 & _will_busy_T_5[31]) begin // @[Rename.scala 70:101]
      map_table_31 <= io_rename_info_bits_1_des_rob;
    end else if (_will_busy_T_1 & _will_busy_T[31]) begin // @[Rename.scala 70:101]
      map_table_31 <= io_rename_info_bits_0_des_rob;
    end
    if (reset) begin // @[Rename.scala 101:23]
      rob_init_info_0_is_valid <= 1'h0; // @[Rename.scala 31:14]
    end else if (io_need_flush) begin // @[Rename.scala 96:22]
      rob_init_info_0_is_valid <= 1'h0; // @[Rename.scala 31:14]
    end else begin
      rob_init_info_0_is_valid <= io_rename_info_bits_0_is_valid; // @[Rename.scala 92:30]
    end
    if (reset) begin // @[Rename.scala 101:23]
      rob_init_info_0_des_rob <= 3'h0; // @[Rename.scala 32:13]
    end else if (io_need_flush) begin // @[Rename.scala 96:22]
      rob_init_info_0_des_rob <= 3'h0; // @[Rename.scala 32:13]
    end else begin
      rob_init_info_0_des_rob <= io_rename_info_bits_0_des_rob; // @[Rename.scala 91:29]
    end
    if (reset) begin // @[Rename.scala 101:23]
      rob_init_info_0_op1_rob <= 3'h0; // @[Rename.scala 33:13]
    end else if (io_need_flush) begin // @[Rename.scala 96:22]
      rob_init_info_0_op1_rob <= 3'h0; // @[Rename.scala 33:13]
    end else if (5'h1f == io_rename_info_bits_0_op1_addr) begin // @[Rename.scala 79:30]
      rob_init_info_0_op1_rob <= map_table_31; // @[Rename.scala 79:30]
    end else if (5'h1e == io_rename_info_bits_0_op1_addr) begin // @[Rename.scala 79:30]
      rob_init_info_0_op1_rob <= map_table_30; // @[Rename.scala 79:30]
    end else begin
      rob_init_info_0_op1_rob <= _GEN_93;
    end
    if (reset) begin // @[Rename.scala 101:23]
      rob_init_info_0_op2_rob <= 3'h0; // @[Rename.scala 34:13]
    end else if (io_need_flush) begin // @[Rename.scala 96:22]
      rob_init_info_0_op2_rob <= 3'h0; // @[Rename.scala 34:13]
    end else if (5'h1f == io_rename_info_bits_0_op2_addr) begin // @[Rename.scala 82:30]
      rob_init_info_0_op2_rob <= map_table_31; // @[Rename.scala 82:30]
    end else if (5'h1e == io_rename_info_bits_0_op2_addr) begin // @[Rename.scala 82:30]
      rob_init_info_0_op2_rob <= map_table_30; // @[Rename.scala 82:30]
    end else begin
      rob_init_info_0_op2_rob <= _GEN_125;
    end
    if (reset) begin // @[Rename.scala 101:23]
      rob_init_info_0_op1_regData <= 32'h0; // @[Rename.scala 35:17]
    end else if (io_need_flush) begin // @[Rename.scala 96:22]
      rob_init_info_0_op1_regData <= 32'h0; // @[Rename.scala 35:17]
    end else begin
      rob_init_info_0_op1_regData <= io_reg_read_0_op1_data; // @[Rename.scala 89:34]
    end
    if (reset) begin // @[Rename.scala 101:23]
      rob_init_info_0_op2_regData <= 32'h0; // @[Rename.scala 36:17]
    end else if (io_need_flush) begin // @[Rename.scala 96:22]
      rob_init_info_0_op2_regData <= 32'h0; // @[Rename.scala 36:17]
    end else begin
      rob_init_info_0_op2_regData <= io_reg_read_0_op2_data; // @[Rename.scala 90:34]
    end
    if (reset) begin // @[Rename.scala 101:23]
      rob_init_info_0_op1_in_rob <= 1'h0; // @[Rename.scala 37:16]
    end else if (io_need_flush) begin // @[Rename.scala 96:22]
      rob_init_info_0_op1_in_rob <= 1'h0; // @[Rename.scala 37:16]
    end else begin
      rob_init_info_0_op1_in_rob <= _rob_init_info_0_op1_in_rob_T[0]; // @[Rename.scala 85:32]
    end
    if (reset) begin // @[Rename.scala 101:23]
      rob_init_info_0_op2_in_rob <= 1'h0; // @[Rename.scala 38:16]
    end else if (io_need_flush) begin // @[Rename.scala 96:22]
      rob_init_info_0_op2_in_rob <= 1'h0; // @[Rename.scala 38:16]
    end else begin
      rob_init_info_0_op2_in_rob <= _rob_init_info_0_op2_in_rob_T[0]; // @[Rename.scala 86:32]
    end
    if (reset) begin // @[Rename.scala 101:23]
      rob_init_info_1_is_valid <= 1'h0; // @[Rename.scala 31:14]
    end else if (io_need_flush) begin // @[Rename.scala 96:22]
      rob_init_info_1_is_valid <= 1'h0; // @[Rename.scala 31:14]
    end else begin
      rob_init_info_1_is_valid <= io_rename_info_bits_1_is_valid; // @[Rename.scala 92:30]
    end
    if (reset) begin // @[Rename.scala 101:23]
      rob_init_info_1_des_rob <= 3'h0; // @[Rename.scala 32:13]
    end else if (io_need_flush) begin // @[Rename.scala 96:22]
      rob_init_info_1_des_rob <= 3'h0; // @[Rename.scala 32:13]
    end else begin
      rob_init_info_1_des_rob <= io_rename_info_bits_1_des_rob; // @[Rename.scala 91:29]
    end
    if (reset) begin // @[Rename.scala 101:23]
      rob_init_info_1_op1_rob <= 3'h0; // @[Rename.scala 33:13]
    end else if (io_need_flush) begin // @[Rename.scala 96:22]
      rob_init_info_1_op1_rob <= 3'h0; // @[Rename.scala 33:13]
    end else if (io_rename_info_bits_0_is_valid & io_rename_info_bits_0_des_addr == io_rename_info_bits_1_op1_addr
      ) begin // @[Rename.scala 80:20]
      rob_init_info_1_op1_rob <= io_rename_info_bits_0_des_rob;
    end else if (5'h1f == io_rename_info_bits_1_op1_addr) begin // @[Rename.scala 80:20]
      rob_init_info_1_op1_rob <= map_table_31; // @[Rename.scala 80:20]
    end else begin
      rob_init_info_1_op1_rob <= _GEN_158;
    end
    if (reset) begin // @[Rename.scala 101:23]
      rob_init_info_1_op2_rob <= 3'h0; // @[Rename.scala 34:13]
    end else if (io_need_flush) begin // @[Rename.scala 96:22]
      rob_init_info_1_op2_rob <= 3'h0; // @[Rename.scala 34:13]
    end else if (io_rename_info_bits_0_is_valid & io_rename_info_bits_0_des_addr == io_rename_info_bits_1_op2_addr
      ) begin // @[Rename.scala 83:20]
      rob_init_info_1_op2_rob <= io_rename_info_bits_0_des_rob;
    end else if (5'h1f == io_rename_info_bits_1_op2_addr) begin // @[Rename.scala 83:20]
      rob_init_info_1_op2_rob <= map_table_31; // @[Rename.scala 83:20]
    end else begin
      rob_init_info_1_op2_rob <= _GEN_190;
    end
    if (reset) begin // @[Rename.scala 101:23]
      rob_init_info_1_op1_regData <= 32'h0; // @[Rename.scala 35:17]
    end else if (io_need_flush) begin // @[Rename.scala 96:22]
      rob_init_info_1_op1_regData <= 32'h0; // @[Rename.scala 35:17]
    end else begin
      rob_init_info_1_op1_regData <= io_reg_read_1_op1_data; // @[Rename.scala 89:34]
    end
    if (reset) begin // @[Rename.scala 101:23]
      rob_init_info_1_op2_regData <= 32'h0; // @[Rename.scala 36:17]
    end else if (io_need_flush) begin // @[Rename.scala 96:22]
      rob_init_info_1_op2_regData <= 32'h0; // @[Rename.scala 36:17]
    end else begin
      rob_init_info_1_op2_regData <= io_reg_read_1_op2_data; // @[Rename.scala 90:34]
    end
    if (reset) begin // @[Rename.scala 101:23]
      rob_init_info_1_op1_in_rob <= 1'h0; // @[Rename.scala 37:16]
    end else if (io_need_flush) begin // @[Rename.scala 96:22]
      rob_init_info_1_op1_in_rob <= 1'h0; // @[Rename.scala 37:16]
    end else begin
      rob_init_info_1_op1_in_rob <= _rob_init_info_1_op1_in_rob_T_4[0] | _rob_init_info_1_op1_rob_T_1 &
        io_rename_info_bits_0_des_addr != 5'h0; // @[Rename.scala 85:32]
    end
    if (reset) begin // @[Rename.scala 101:23]
      rob_init_info_1_op2_in_rob <= 1'h0; // @[Rename.scala 38:16]
    end else if (io_need_flush) begin // @[Rename.scala 96:22]
      rob_init_info_1_op2_in_rob <= 1'h0; // @[Rename.scala 38:16]
    end else begin
      rob_init_info_1_op2_in_rob <= _rob_init_info_1_op2_in_rob_T_4[0] | _rob_init_info_1_op2_rob_T_1 &
        _rob_init_info_1_op1_in_rob_T_2; // @[Rename.scala 86:32]
    end
    if (reset) begin // @[Rename.scala 74:36]
      rob_init_info_valid <= 1'h0; // @[Rename.scala 74:36]
    end else if (io_need_flush) begin // @[Rename.scala 96:22]
      rob_init_info_valid <= 1'h0; // @[Rename.scala 98:24]
    end else begin
      rob_init_info_valid <= io_rename_info_valid; // @[Rename.scala 94:22]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  busy_table = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  map_table_1 = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  map_table_2 = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  map_table_3 = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  map_table_4 = _RAND_4[2:0];
  _RAND_5 = {1{`RANDOM}};
  map_table_5 = _RAND_5[2:0];
  _RAND_6 = {1{`RANDOM}};
  map_table_6 = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  map_table_7 = _RAND_7[2:0];
  _RAND_8 = {1{`RANDOM}};
  map_table_8 = _RAND_8[2:0];
  _RAND_9 = {1{`RANDOM}};
  map_table_9 = _RAND_9[2:0];
  _RAND_10 = {1{`RANDOM}};
  map_table_10 = _RAND_10[2:0];
  _RAND_11 = {1{`RANDOM}};
  map_table_11 = _RAND_11[2:0];
  _RAND_12 = {1{`RANDOM}};
  map_table_12 = _RAND_12[2:0];
  _RAND_13 = {1{`RANDOM}};
  map_table_13 = _RAND_13[2:0];
  _RAND_14 = {1{`RANDOM}};
  map_table_14 = _RAND_14[2:0];
  _RAND_15 = {1{`RANDOM}};
  map_table_15 = _RAND_15[2:0];
  _RAND_16 = {1{`RANDOM}};
  map_table_16 = _RAND_16[2:0];
  _RAND_17 = {1{`RANDOM}};
  map_table_17 = _RAND_17[2:0];
  _RAND_18 = {1{`RANDOM}};
  map_table_18 = _RAND_18[2:0];
  _RAND_19 = {1{`RANDOM}};
  map_table_19 = _RAND_19[2:0];
  _RAND_20 = {1{`RANDOM}};
  map_table_20 = _RAND_20[2:0];
  _RAND_21 = {1{`RANDOM}};
  map_table_21 = _RAND_21[2:0];
  _RAND_22 = {1{`RANDOM}};
  map_table_22 = _RAND_22[2:0];
  _RAND_23 = {1{`RANDOM}};
  map_table_23 = _RAND_23[2:0];
  _RAND_24 = {1{`RANDOM}};
  map_table_24 = _RAND_24[2:0];
  _RAND_25 = {1{`RANDOM}};
  map_table_25 = _RAND_25[2:0];
  _RAND_26 = {1{`RANDOM}};
  map_table_26 = _RAND_26[2:0];
  _RAND_27 = {1{`RANDOM}};
  map_table_27 = _RAND_27[2:0];
  _RAND_28 = {1{`RANDOM}};
  map_table_28 = _RAND_28[2:0];
  _RAND_29 = {1{`RANDOM}};
  map_table_29 = _RAND_29[2:0];
  _RAND_30 = {1{`RANDOM}};
  map_table_30 = _RAND_30[2:0];
  _RAND_31 = {1{`RANDOM}};
  map_table_31 = _RAND_31[2:0];
  _RAND_32 = {1{`RANDOM}};
  rob_init_info_0_is_valid = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  rob_init_info_0_des_rob = _RAND_33[2:0];
  _RAND_34 = {1{`RANDOM}};
  rob_init_info_0_op1_rob = _RAND_34[2:0];
  _RAND_35 = {1{`RANDOM}};
  rob_init_info_0_op2_rob = _RAND_35[2:0];
  _RAND_36 = {1{`RANDOM}};
  rob_init_info_0_op1_regData = _RAND_36[31:0];
  _RAND_37 = {1{`RANDOM}};
  rob_init_info_0_op2_regData = _RAND_37[31:0];
  _RAND_38 = {1{`RANDOM}};
  rob_init_info_0_op1_in_rob = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  rob_init_info_0_op2_in_rob = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  rob_init_info_1_is_valid = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  rob_init_info_1_des_rob = _RAND_41[2:0];
  _RAND_42 = {1{`RANDOM}};
  rob_init_info_1_op1_rob = _RAND_42[2:0];
  _RAND_43 = {1{`RANDOM}};
  rob_init_info_1_op2_rob = _RAND_43[2:0];
  _RAND_44 = {1{`RANDOM}};
  rob_init_info_1_op1_regData = _RAND_44[31:0];
  _RAND_45 = {1{`RANDOM}};
  rob_init_info_1_op2_regData = _RAND_45[31:0];
  _RAND_46 = {1{`RANDOM}};
  rob_init_info_1_op1_in_rob = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  rob_init_info_1_op2_in_rob = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  rob_init_info_valid = _RAND_48[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Regfile(
  input         clock,
  input         reset,
  input  [4:0]  io_reg_read_0_op1_addr,
  input  [4:0]  io_reg_read_0_op2_addr,
  output [31:0] io_reg_read_0_op1_data,
  output [31:0] io_reg_read_0_op2_data,
  input  [4:0]  io_reg_read_1_op1_addr,
  input  [4:0]  io_reg_read_1_op2_addr,
  output [31:0] io_reg_read_1_op1_data,
  output [31:0] io_reg_read_1_op2_data,
  input         io_rob_commit_i_0_valid,
  input  [4:0]  io_rob_commit_i_0_bits_commit_addr,
  input  [31:0] io_rob_commit_i_0_bits_commit_data,
  input         io_rob_commit_i_1_valid,
  input  [4:0]  io_rob_commit_i_1_bits_commit_addr,
  input  [31:0] io_rob_commit_i_1_bits_commit_data
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] regfile_1; // @[Regfile.scala 18:24]
  reg [31:0] regfile_2; // @[Regfile.scala 18:24]
  reg [31:0] regfile_3; // @[Regfile.scala 18:24]
  reg [31:0] regfile_4; // @[Regfile.scala 18:24]
  reg [31:0] regfile_5; // @[Regfile.scala 18:24]
  reg [31:0] regfile_6; // @[Regfile.scala 18:24]
  reg [31:0] regfile_7; // @[Regfile.scala 18:24]
  reg [31:0] regfile_8; // @[Regfile.scala 18:24]
  reg [31:0] regfile_9; // @[Regfile.scala 18:24]
  reg [31:0] regfile_10; // @[Regfile.scala 18:24]
  reg [31:0] regfile_11; // @[Regfile.scala 18:24]
  reg [31:0] regfile_12; // @[Regfile.scala 18:24]
  reg [31:0] regfile_13; // @[Regfile.scala 18:24]
  reg [31:0] regfile_14; // @[Regfile.scala 18:24]
  reg [31:0] regfile_15; // @[Regfile.scala 18:24]
  reg [31:0] regfile_16; // @[Regfile.scala 18:24]
  reg [31:0] regfile_17; // @[Regfile.scala 18:24]
  reg [31:0] regfile_18; // @[Regfile.scala 18:24]
  reg [31:0] regfile_19; // @[Regfile.scala 18:24]
  reg [31:0] regfile_20; // @[Regfile.scala 18:24]
  reg [31:0] regfile_21; // @[Regfile.scala 18:24]
  reg [31:0] regfile_22; // @[Regfile.scala 18:24]
  reg [31:0] regfile_23; // @[Regfile.scala 18:24]
  reg [31:0] regfile_24; // @[Regfile.scala 18:24]
  reg [31:0] regfile_25; // @[Regfile.scala 18:24]
  reg [31:0] regfile_26; // @[Regfile.scala 18:24]
  reg [31:0] regfile_27; // @[Regfile.scala 18:24]
  reg [31:0] regfile_28; // @[Regfile.scala 18:24]
  reg [31:0] regfile_29; // @[Regfile.scala 18:24]
  reg [31:0] regfile_30; // @[Regfile.scala 18:24]
  reg [31:0] regfile_31; // @[Regfile.scala 18:24]
  wire [31:0] commit_idx_0 = 32'h1 << io_rob_commit_i_0_bits_commit_addr; // @[OneHot.scala 58:35]
  wire [31:0] commit_idx_1 = 32'h1 << io_rob_commit_i_1_bits_commit_addr; // @[OneHot.scala 58:35]
  wire [31:0] _next_data_1_T_2 = io_rob_commit_i_0_valid & commit_idx_0[1] ? io_rob_commit_i_0_bits_commit_data :
    regfile_1; // @[Regfile.scala 25:93]
  wire [31:0] next_data_1 = io_rob_commit_i_1_valid & commit_idx_1[1] ? io_rob_commit_i_1_bits_commit_data :
    _next_data_1_T_2; // @[Regfile.scala 25:93]
  wire [31:0] _next_data_2_T_2 = io_rob_commit_i_0_valid & commit_idx_0[2] ? io_rob_commit_i_0_bits_commit_data :
    regfile_2; // @[Regfile.scala 25:93]
  wire [31:0] next_data_2 = io_rob_commit_i_1_valid & commit_idx_1[2] ? io_rob_commit_i_1_bits_commit_data :
    _next_data_2_T_2; // @[Regfile.scala 25:93]
  wire [31:0] _next_data_3_T_2 = io_rob_commit_i_0_valid & commit_idx_0[3] ? io_rob_commit_i_0_bits_commit_data :
    regfile_3; // @[Regfile.scala 25:93]
  wire [31:0] next_data_3 = io_rob_commit_i_1_valid & commit_idx_1[3] ? io_rob_commit_i_1_bits_commit_data :
    _next_data_3_T_2; // @[Regfile.scala 25:93]
  wire [31:0] _next_data_4_T_2 = io_rob_commit_i_0_valid & commit_idx_0[4] ? io_rob_commit_i_0_bits_commit_data :
    regfile_4; // @[Regfile.scala 25:93]
  wire [31:0] next_data_4 = io_rob_commit_i_1_valid & commit_idx_1[4] ? io_rob_commit_i_1_bits_commit_data :
    _next_data_4_T_2; // @[Regfile.scala 25:93]
  wire [31:0] _next_data_5_T_2 = io_rob_commit_i_0_valid & commit_idx_0[5] ? io_rob_commit_i_0_bits_commit_data :
    regfile_5; // @[Regfile.scala 25:93]
  wire [31:0] next_data_5 = io_rob_commit_i_1_valid & commit_idx_1[5] ? io_rob_commit_i_1_bits_commit_data :
    _next_data_5_T_2; // @[Regfile.scala 25:93]
  wire [31:0] _next_data_6_T_2 = io_rob_commit_i_0_valid & commit_idx_0[6] ? io_rob_commit_i_0_bits_commit_data :
    regfile_6; // @[Regfile.scala 25:93]
  wire [31:0] next_data_6 = io_rob_commit_i_1_valid & commit_idx_1[6] ? io_rob_commit_i_1_bits_commit_data :
    _next_data_6_T_2; // @[Regfile.scala 25:93]
  wire [31:0] _next_data_7_T_2 = io_rob_commit_i_0_valid & commit_idx_0[7] ? io_rob_commit_i_0_bits_commit_data :
    regfile_7; // @[Regfile.scala 25:93]
  wire [31:0] next_data_7 = io_rob_commit_i_1_valid & commit_idx_1[7] ? io_rob_commit_i_1_bits_commit_data :
    _next_data_7_T_2; // @[Regfile.scala 25:93]
  wire [31:0] _next_data_8_T_2 = io_rob_commit_i_0_valid & commit_idx_0[8] ? io_rob_commit_i_0_bits_commit_data :
    regfile_8; // @[Regfile.scala 25:93]
  wire [31:0] next_data_8 = io_rob_commit_i_1_valid & commit_idx_1[8] ? io_rob_commit_i_1_bits_commit_data :
    _next_data_8_T_2; // @[Regfile.scala 25:93]
  wire [31:0] _next_data_9_T_2 = io_rob_commit_i_0_valid & commit_idx_0[9] ? io_rob_commit_i_0_bits_commit_data :
    regfile_9; // @[Regfile.scala 25:93]
  wire [31:0] next_data_9 = io_rob_commit_i_1_valid & commit_idx_1[9] ? io_rob_commit_i_1_bits_commit_data :
    _next_data_9_T_2; // @[Regfile.scala 25:93]
  wire [31:0] _next_data_10_T_2 = io_rob_commit_i_0_valid & commit_idx_0[10] ? io_rob_commit_i_0_bits_commit_data :
    regfile_10; // @[Regfile.scala 25:93]
  wire [31:0] next_data_10 = io_rob_commit_i_1_valid & commit_idx_1[10] ? io_rob_commit_i_1_bits_commit_data :
    _next_data_10_T_2; // @[Regfile.scala 25:93]
  wire [31:0] _next_data_11_T_2 = io_rob_commit_i_0_valid & commit_idx_0[11] ? io_rob_commit_i_0_bits_commit_data :
    regfile_11; // @[Regfile.scala 25:93]
  wire [31:0] next_data_11 = io_rob_commit_i_1_valid & commit_idx_1[11] ? io_rob_commit_i_1_bits_commit_data :
    _next_data_11_T_2; // @[Regfile.scala 25:93]
  wire [31:0] _next_data_12_T_2 = io_rob_commit_i_0_valid & commit_idx_0[12] ? io_rob_commit_i_0_bits_commit_data :
    regfile_12; // @[Regfile.scala 25:93]
  wire [31:0] next_data_12 = io_rob_commit_i_1_valid & commit_idx_1[12] ? io_rob_commit_i_1_bits_commit_data :
    _next_data_12_T_2; // @[Regfile.scala 25:93]
  wire [31:0] _next_data_13_T_2 = io_rob_commit_i_0_valid & commit_idx_0[13] ? io_rob_commit_i_0_bits_commit_data :
    regfile_13; // @[Regfile.scala 25:93]
  wire [31:0] next_data_13 = io_rob_commit_i_1_valid & commit_idx_1[13] ? io_rob_commit_i_1_bits_commit_data :
    _next_data_13_T_2; // @[Regfile.scala 25:93]
  wire [31:0] _next_data_14_T_2 = io_rob_commit_i_0_valid & commit_idx_0[14] ? io_rob_commit_i_0_bits_commit_data :
    regfile_14; // @[Regfile.scala 25:93]
  wire [31:0] next_data_14 = io_rob_commit_i_1_valid & commit_idx_1[14] ? io_rob_commit_i_1_bits_commit_data :
    _next_data_14_T_2; // @[Regfile.scala 25:93]
  wire [31:0] _next_data_15_T_2 = io_rob_commit_i_0_valid & commit_idx_0[15] ? io_rob_commit_i_0_bits_commit_data :
    regfile_15; // @[Regfile.scala 25:93]
  wire [31:0] next_data_15 = io_rob_commit_i_1_valid & commit_idx_1[15] ? io_rob_commit_i_1_bits_commit_data :
    _next_data_15_T_2; // @[Regfile.scala 25:93]
  wire [31:0] _next_data_16_T_2 = io_rob_commit_i_0_valid & commit_idx_0[16] ? io_rob_commit_i_0_bits_commit_data :
    regfile_16; // @[Regfile.scala 25:93]
  wire [31:0] next_data_16 = io_rob_commit_i_1_valid & commit_idx_1[16] ? io_rob_commit_i_1_bits_commit_data :
    _next_data_16_T_2; // @[Regfile.scala 25:93]
  wire [31:0] _next_data_17_T_2 = io_rob_commit_i_0_valid & commit_idx_0[17] ? io_rob_commit_i_0_bits_commit_data :
    regfile_17; // @[Regfile.scala 25:93]
  wire [31:0] next_data_17 = io_rob_commit_i_1_valid & commit_idx_1[17] ? io_rob_commit_i_1_bits_commit_data :
    _next_data_17_T_2; // @[Regfile.scala 25:93]
  wire [31:0] _next_data_18_T_2 = io_rob_commit_i_0_valid & commit_idx_0[18] ? io_rob_commit_i_0_bits_commit_data :
    regfile_18; // @[Regfile.scala 25:93]
  wire [31:0] next_data_18 = io_rob_commit_i_1_valid & commit_idx_1[18] ? io_rob_commit_i_1_bits_commit_data :
    _next_data_18_T_2; // @[Regfile.scala 25:93]
  wire [31:0] _next_data_19_T_2 = io_rob_commit_i_0_valid & commit_idx_0[19] ? io_rob_commit_i_0_bits_commit_data :
    regfile_19; // @[Regfile.scala 25:93]
  wire [31:0] next_data_19 = io_rob_commit_i_1_valid & commit_idx_1[19] ? io_rob_commit_i_1_bits_commit_data :
    _next_data_19_T_2; // @[Regfile.scala 25:93]
  wire [31:0] _next_data_20_T_2 = io_rob_commit_i_0_valid & commit_idx_0[20] ? io_rob_commit_i_0_bits_commit_data :
    regfile_20; // @[Regfile.scala 25:93]
  wire [31:0] next_data_20 = io_rob_commit_i_1_valid & commit_idx_1[20] ? io_rob_commit_i_1_bits_commit_data :
    _next_data_20_T_2; // @[Regfile.scala 25:93]
  wire [31:0] _next_data_21_T_2 = io_rob_commit_i_0_valid & commit_idx_0[21] ? io_rob_commit_i_0_bits_commit_data :
    regfile_21; // @[Regfile.scala 25:93]
  wire [31:0] next_data_21 = io_rob_commit_i_1_valid & commit_idx_1[21] ? io_rob_commit_i_1_bits_commit_data :
    _next_data_21_T_2; // @[Regfile.scala 25:93]
  wire [31:0] _next_data_22_T_2 = io_rob_commit_i_0_valid & commit_idx_0[22] ? io_rob_commit_i_0_bits_commit_data :
    regfile_22; // @[Regfile.scala 25:93]
  wire [31:0] next_data_22 = io_rob_commit_i_1_valid & commit_idx_1[22] ? io_rob_commit_i_1_bits_commit_data :
    _next_data_22_T_2; // @[Regfile.scala 25:93]
  wire [31:0] _next_data_23_T_2 = io_rob_commit_i_0_valid & commit_idx_0[23] ? io_rob_commit_i_0_bits_commit_data :
    regfile_23; // @[Regfile.scala 25:93]
  wire [31:0] next_data_23 = io_rob_commit_i_1_valid & commit_idx_1[23] ? io_rob_commit_i_1_bits_commit_data :
    _next_data_23_T_2; // @[Regfile.scala 25:93]
  wire [31:0] _next_data_24_T_2 = io_rob_commit_i_0_valid & commit_idx_0[24] ? io_rob_commit_i_0_bits_commit_data :
    regfile_24; // @[Regfile.scala 25:93]
  wire [31:0] next_data_24 = io_rob_commit_i_1_valid & commit_idx_1[24] ? io_rob_commit_i_1_bits_commit_data :
    _next_data_24_T_2; // @[Regfile.scala 25:93]
  wire [31:0] _next_data_25_T_2 = io_rob_commit_i_0_valid & commit_idx_0[25] ? io_rob_commit_i_0_bits_commit_data :
    regfile_25; // @[Regfile.scala 25:93]
  wire [31:0] next_data_25 = io_rob_commit_i_1_valid & commit_idx_1[25] ? io_rob_commit_i_1_bits_commit_data :
    _next_data_25_T_2; // @[Regfile.scala 25:93]
  wire [31:0] _next_data_26_T_2 = io_rob_commit_i_0_valid & commit_idx_0[26] ? io_rob_commit_i_0_bits_commit_data :
    regfile_26; // @[Regfile.scala 25:93]
  wire [31:0] next_data_26 = io_rob_commit_i_1_valid & commit_idx_1[26] ? io_rob_commit_i_1_bits_commit_data :
    _next_data_26_T_2; // @[Regfile.scala 25:93]
  wire [31:0] _next_data_27_T_2 = io_rob_commit_i_0_valid & commit_idx_0[27] ? io_rob_commit_i_0_bits_commit_data :
    regfile_27; // @[Regfile.scala 25:93]
  wire [31:0] next_data_27 = io_rob_commit_i_1_valid & commit_idx_1[27] ? io_rob_commit_i_1_bits_commit_data :
    _next_data_27_T_2; // @[Regfile.scala 25:93]
  wire [31:0] _next_data_28_T_2 = io_rob_commit_i_0_valid & commit_idx_0[28] ? io_rob_commit_i_0_bits_commit_data :
    regfile_28; // @[Regfile.scala 25:93]
  wire [31:0] next_data_28 = io_rob_commit_i_1_valid & commit_idx_1[28] ? io_rob_commit_i_1_bits_commit_data :
    _next_data_28_T_2; // @[Regfile.scala 25:93]
  wire [31:0] _next_data_29_T_2 = io_rob_commit_i_0_valid & commit_idx_0[29] ? io_rob_commit_i_0_bits_commit_data :
    regfile_29; // @[Regfile.scala 25:93]
  wire [31:0] next_data_29 = io_rob_commit_i_1_valid & commit_idx_1[29] ? io_rob_commit_i_1_bits_commit_data :
    _next_data_29_T_2; // @[Regfile.scala 25:93]
  wire [31:0] _next_data_30_T_2 = io_rob_commit_i_0_valid & commit_idx_0[30] ? io_rob_commit_i_0_bits_commit_data :
    regfile_30; // @[Regfile.scala 25:93]
  wire [31:0] next_data_30 = io_rob_commit_i_1_valid & commit_idx_1[30] ? io_rob_commit_i_1_bits_commit_data :
    _next_data_30_T_2; // @[Regfile.scala 25:93]
  wire [31:0] _next_data_31_T_2 = io_rob_commit_i_0_valid & commit_idx_0[31] ? io_rob_commit_i_0_bits_commit_data :
    regfile_31; // @[Regfile.scala 25:93]
  wire [31:0] next_data_31 = io_rob_commit_i_1_valid & commit_idx_1[31] ? io_rob_commit_i_1_bits_commit_data :
    _next_data_31_T_2; // @[Regfile.scala 25:93]
  wire [31:0] _GEN_1 = 5'h1 == io_reg_read_0_op1_addr ? next_data_1 : 32'h0; // @[Regfile.scala 29:28 Regfile.scala 29:28]
  wire [31:0] _GEN_2 = 5'h2 == io_reg_read_0_op1_addr ? next_data_2 : _GEN_1; // @[Regfile.scala 29:28 Regfile.scala 29:28]
  wire [31:0] _GEN_3 = 5'h3 == io_reg_read_0_op1_addr ? next_data_3 : _GEN_2; // @[Regfile.scala 29:28 Regfile.scala 29:28]
  wire [31:0] _GEN_4 = 5'h4 == io_reg_read_0_op1_addr ? next_data_4 : _GEN_3; // @[Regfile.scala 29:28 Regfile.scala 29:28]
  wire [31:0] _GEN_5 = 5'h5 == io_reg_read_0_op1_addr ? next_data_5 : _GEN_4; // @[Regfile.scala 29:28 Regfile.scala 29:28]
  wire [31:0] _GEN_6 = 5'h6 == io_reg_read_0_op1_addr ? next_data_6 : _GEN_5; // @[Regfile.scala 29:28 Regfile.scala 29:28]
  wire [31:0] _GEN_7 = 5'h7 == io_reg_read_0_op1_addr ? next_data_7 : _GEN_6; // @[Regfile.scala 29:28 Regfile.scala 29:28]
  wire [31:0] _GEN_8 = 5'h8 == io_reg_read_0_op1_addr ? next_data_8 : _GEN_7; // @[Regfile.scala 29:28 Regfile.scala 29:28]
  wire [31:0] _GEN_9 = 5'h9 == io_reg_read_0_op1_addr ? next_data_9 : _GEN_8; // @[Regfile.scala 29:28 Regfile.scala 29:28]
  wire [31:0] _GEN_10 = 5'ha == io_reg_read_0_op1_addr ? next_data_10 : _GEN_9; // @[Regfile.scala 29:28 Regfile.scala 29:28]
  wire [31:0] _GEN_11 = 5'hb == io_reg_read_0_op1_addr ? next_data_11 : _GEN_10; // @[Regfile.scala 29:28 Regfile.scala 29:28]
  wire [31:0] _GEN_12 = 5'hc == io_reg_read_0_op1_addr ? next_data_12 : _GEN_11; // @[Regfile.scala 29:28 Regfile.scala 29:28]
  wire [31:0] _GEN_13 = 5'hd == io_reg_read_0_op1_addr ? next_data_13 : _GEN_12; // @[Regfile.scala 29:28 Regfile.scala 29:28]
  wire [31:0] _GEN_14 = 5'he == io_reg_read_0_op1_addr ? next_data_14 : _GEN_13; // @[Regfile.scala 29:28 Regfile.scala 29:28]
  wire [31:0] _GEN_15 = 5'hf == io_reg_read_0_op1_addr ? next_data_15 : _GEN_14; // @[Regfile.scala 29:28 Regfile.scala 29:28]
  wire [31:0] _GEN_16 = 5'h10 == io_reg_read_0_op1_addr ? next_data_16 : _GEN_15; // @[Regfile.scala 29:28 Regfile.scala 29:28]
  wire [31:0] _GEN_17 = 5'h11 == io_reg_read_0_op1_addr ? next_data_17 : _GEN_16; // @[Regfile.scala 29:28 Regfile.scala 29:28]
  wire [31:0] _GEN_18 = 5'h12 == io_reg_read_0_op1_addr ? next_data_18 : _GEN_17; // @[Regfile.scala 29:28 Regfile.scala 29:28]
  wire [31:0] _GEN_19 = 5'h13 == io_reg_read_0_op1_addr ? next_data_19 : _GEN_18; // @[Regfile.scala 29:28 Regfile.scala 29:28]
  wire [31:0] _GEN_20 = 5'h14 == io_reg_read_0_op1_addr ? next_data_20 : _GEN_19; // @[Regfile.scala 29:28 Regfile.scala 29:28]
  wire [31:0] _GEN_21 = 5'h15 == io_reg_read_0_op1_addr ? next_data_21 : _GEN_20; // @[Regfile.scala 29:28 Regfile.scala 29:28]
  wire [31:0] _GEN_22 = 5'h16 == io_reg_read_0_op1_addr ? next_data_22 : _GEN_21; // @[Regfile.scala 29:28 Regfile.scala 29:28]
  wire [31:0] _GEN_23 = 5'h17 == io_reg_read_0_op1_addr ? next_data_23 : _GEN_22; // @[Regfile.scala 29:28 Regfile.scala 29:28]
  wire [31:0] _GEN_24 = 5'h18 == io_reg_read_0_op1_addr ? next_data_24 : _GEN_23; // @[Regfile.scala 29:28 Regfile.scala 29:28]
  wire [31:0] _GEN_25 = 5'h19 == io_reg_read_0_op1_addr ? next_data_25 : _GEN_24; // @[Regfile.scala 29:28 Regfile.scala 29:28]
  wire [31:0] _GEN_26 = 5'h1a == io_reg_read_0_op1_addr ? next_data_26 : _GEN_25; // @[Regfile.scala 29:28 Regfile.scala 29:28]
  wire [31:0] _GEN_27 = 5'h1b == io_reg_read_0_op1_addr ? next_data_27 : _GEN_26; // @[Regfile.scala 29:28 Regfile.scala 29:28]
  wire [31:0] _GEN_28 = 5'h1c == io_reg_read_0_op1_addr ? next_data_28 : _GEN_27; // @[Regfile.scala 29:28 Regfile.scala 29:28]
  wire [31:0] _GEN_29 = 5'h1d == io_reg_read_0_op1_addr ? next_data_29 : _GEN_28; // @[Regfile.scala 29:28 Regfile.scala 29:28]
  wire [31:0] _GEN_30 = 5'h1e == io_reg_read_0_op1_addr ? next_data_30 : _GEN_29; // @[Regfile.scala 29:28 Regfile.scala 29:28]
  wire [31:0] _GEN_33 = 5'h1 == io_reg_read_0_op2_addr ? next_data_1 : 32'h0; // @[Regfile.scala 30:28 Regfile.scala 30:28]
  wire [31:0] _GEN_34 = 5'h2 == io_reg_read_0_op2_addr ? next_data_2 : _GEN_33; // @[Regfile.scala 30:28 Regfile.scala 30:28]
  wire [31:0] _GEN_35 = 5'h3 == io_reg_read_0_op2_addr ? next_data_3 : _GEN_34; // @[Regfile.scala 30:28 Regfile.scala 30:28]
  wire [31:0] _GEN_36 = 5'h4 == io_reg_read_0_op2_addr ? next_data_4 : _GEN_35; // @[Regfile.scala 30:28 Regfile.scala 30:28]
  wire [31:0] _GEN_37 = 5'h5 == io_reg_read_0_op2_addr ? next_data_5 : _GEN_36; // @[Regfile.scala 30:28 Regfile.scala 30:28]
  wire [31:0] _GEN_38 = 5'h6 == io_reg_read_0_op2_addr ? next_data_6 : _GEN_37; // @[Regfile.scala 30:28 Regfile.scala 30:28]
  wire [31:0] _GEN_39 = 5'h7 == io_reg_read_0_op2_addr ? next_data_7 : _GEN_38; // @[Regfile.scala 30:28 Regfile.scala 30:28]
  wire [31:0] _GEN_40 = 5'h8 == io_reg_read_0_op2_addr ? next_data_8 : _GEN_39; // @[Regfile.scala 30:28 Regfile.scala 30:28]
  wire [31:0] _GEN_41 = 5'h9 == io_reg_read_0_op2_addr ? next_data_9 : _GEN_40; // @[Regfile.scala 30:28 Regfile.scala 30:28]
  wire [31:0] _GEN_42 = 5'ha == io_reg_read_0_op2_addr ? next_data_10 : _GEN_41; // @[Regfile.scala 30:28 Regfile.scala 30:28]
  wire [31:0] _GEN_43 = 5'hb == io_reg_read_0_op2_addr ? next_data_11 : _GEN_42; // @[Regfile.scala 30:28 Regfile.scala 30:28]
  wire [31:0] _GEN_44 = 5'hc == io_reg_read_0_op2_addr ? next_data_12 : _GEN_43; // @[Regfile.scala 30:28 Regfile.scala 30:28]
  wire [31:0] _GEN_45 = 5'hd == io_reg_read_0_op2_addr ? next_data_13 : _GEN_44; // @[Regfile.scala 30:28 Regfile.scala 30:28]
  wire [31:0] _GEN_46 = 5'he == io_reg_read_0_op2_addr ? next_data_14 : _GEN_45; // @[Regfile.scala 30:28 Regfile.scala 30:28]
  wire [31:0] _GEN_47 = 5'hf == io_reg_read_0_op2_addr ? next_data_15 : _GEN_46; // @[Regfile.scala 30:28 Regfile.scala 30:28]
  wire [31:0] _GEN_48 = 5'h10 == io_reg_read_0_op2_addr ? next_data_16 : _GEN_47; // @[Regfile.scala 30:28 Regfile.scala 30:28]
  wire [31:0] _GEN_49 = 5'h11 == io_reg_read_0_op2_addr ? next_data_17 : _GEN_48; // @[Regfile.scala 30:28 Regfile.scala 30:28]
  wire [31:0] _GEN_50 = 5'h12 == io_reg_read_0_op2_addr ? next_data_18 : _GEN_49; // @[Regfile.scala 30:28 Regfile.scala 30:28]
  wire [31:0] _GEN_51 = 5'h13 == io_reg_read_0_op2_addr ? next_data_19 : _GEN_50; // @[Regfile.scala 30:28 Regfile.scala 30:28]
  wire [31:0] _GEN_52 = 5'h14 == io_reg_read_0_op2_addr ? next_data_20 : _GEN_51; // @[Regfile.scala 30:28 Regfile.scala 30:28]
  wire [31:0] _GEN_53 = 5'h15 == io_reg_read_0_op2_addr ? next_data_21 : _GEN_52; // @[Regfile.scala 30:28 Regfile.scala 30:28]
  wire [31:0] _GEN_54 = 5'h16 == io_reg_read_0_op2_addr ? next_data_22 : _GEN_53; // @[Regfile.scala 30:28 Regfile.scala 30:28]
  wire [31:0] _GEN_55 = 5'h17 == io_reg_read_0_op2_addr ? next_data_23 : _GEN_54; // @[Regfile.scala 30:28 Regfile.scala 30:28]
  wire [31:0] _GEN_56 = 5'h18 == io_reg_read_0_op2_addr ? next_data_24 : _GEN_55; // @[Regfile.scala 30:28 Regfile.scala 30:28]
  wire [31:0] _GEN_57 = 5'h19 == io_reg_read_0_op2_addr ? next_data_25 : _GEN_56; // @[Regfile.scala 30:28 Regfile.scala 30:28]
  wire [31:0] _GEN_58 = 5'h1a == io_reg_read_0_op2_addr ? next_data_26 : _GEN_57; // @[Regfile.scala 30:28 Regfile.scala 30:28]
  wire [31:0] _GEN_59 = 5'h1b == io_reg_read_0_op2_addr ? next_data_27 : _GEN_58; // @[Regfile.scala 30:28 Regfile.scala 30:28]
  wire [31:0] _GEN_60 = 5'h1c == io_reg_read_0_op2_addr ? next_data_28 : _GEN_59; // @[Regfile.scala 30:28 Regfile.scala 30:28]
  wire [31:0] _GEN_61 = 5'h1d == io_reg_read_0_op2_addr ? next_data_29 : _GEN_60; // @[Regfile.scala 30:28 Regfile.scala 30:28]
  wire [31:0] _GEN_62 = 5'h1e == io_reg_read_0_op2_addr ? next_data_30 : _GEN_61; // @[Regfile.scala 30:28 Regfile.scala 30:28]
  wire [31:0] _GEN_65 = 5'h1 == io_reg_read_1_op1_addr ? next_data_1 : 32'h0; // @[Regfile.scala 29:28 Regfile.scala 29:28]
  wire [31:0] _GEN_66 = 5'h2 == io_reg_read_1_op1_addr ? next_data_2 : _GEN_65; // @[Regfile.scala 29:28 Regfile.scala 29:28]
  wire [31:0] _GEN_67 = 5'h3 == io_reg_read_1_op1_addr ? next_data_3 : _GEN_66; // @[Regfile.scala 29:28 Regfile.scala 29:28]
  wire [31:0] _GEN_68 = 5'h4 == io_reg_read_1_op1_addr ? next_data_4 : _GEN_67; // @[Regfile.scala 29:28 Regfile.scala 29:28]
  wire [31:0] _GEN_69 = 5'h5 == io_reg_read_1_op1_addr ? next_data_5 : _GEN_68; // @[Regfile.scala 29:28 Regfile.scala 29:28]
  wire [31:0] _GEN_70 = 5'h6 == io_reg_read_1_op1_addr ? next_data_6 : _GEN_69; // @[Regfile.scala 29:28 Regfile.scala 29:28]
  wire [31:0] _GEN_71 = 5'h7 == io_reg_read_1_op1_addr ? next_data_7 : _GEN_70; // @[Regfile.scala 29:28 Regfile.scala 29:28]
  wire [31:0] _GEN_72 = 5'h8 == io_reg_read_1_op1_addr ? next_data_8 : _GEN_71; // @[Regfile.scala 29:28 Regfile.scala 29:28]
  wire [31:0] _GEN_73 = 5'h9 == io_reg_read_1_op1_addr ? next_data_9 : _GEN_72; // @[Regfile.scala 29:28 Regfile.scala 29:28]
  wire [31:0] _GEN_74 = 5'ha == io_reg_read_1_op1_addr ? next_data_10 : _GEN_73; // @[Regfile.scala 29:28 Regfile.scala 29:28]
  wire [31:0] _GEN_75 = 5'hb == io_reg_read_1_op1_addr ? next_data_11 : _GEN_74; // @[Regfile.scala 29:28 Regfile.scala 29:28]
  wire [31:0] _GEN_76 = 5'hc == io_reg_read_1_op1_addr ? next_data_12 : _GEN_75; // @[Regfile.scala 29:28 Regfile.scala 29:28]
  wire [31:0] _GEN_77 = 5'hd == io_reg_read_1_op1_addr ? next_data_13 : _GEN_76; // @[Regfile.scala 29:28 Regfile.scala 29:28]
  wire [31:0] _GEN_78 = 5'he == io_reg_read_1_op1_addr ? next_data_14 : _GEN_77; // @[Regfile.scala 29:28 Regfile.scala 29:28]
  wire [31:0] _GEN_79 = 5'hf == io_reg_read_1_op1_addr ? next_data_15 : _GEN_78; // @[Regfile.scala 29:28 Regfile.scala 29:28]
  wire [31:0] _GEN_80 = 5'h10 == io_reg_read_1_op1_addr ? next_data_16 : _GEN_79; // @[Regfile.scala 29:28 Regfile.scala 29:28]
  wire [31:0] _GEN_81 = 5'h11 == io_reg_read_1_op1_addr ? next_data_17 : _GEN_80; // @[Regfile.scala 29:28 Regfile.scala 29:28]
  wire [31:0] _GEN_82 = 5'h12 == io_reg_read_1_op1_addr ? next_data_18 : _GEN_81; // @[Regfile.scala 29:28 Regfile.scala 29:28]
  wire [31:0] _GEN_83 = 5'h13 == io_reg_read_1_op1_addr ? next_data_19 : _GEN_82; // @[Regfile.scala 29:28 Regfile.scala 29:28]
  wire [31:0] _GEN_84 = 5'h14 == io_reg_read_1_op1_addr ? next_data_20 : _GEN_83; // @[Regfile.scala 29:28 Regfile.scala 29:28]
  wire [31:0] _GEN_85 = 5'h15 == io_reg_read_1_op1_addr ? next_data_21 : _GEN_84; // @[Regfile.scala 29:28 Regfile.scala 29:28]
  wire [31:0] _GEN_86 = 5'h16 == io_reg_read_1_op1_addr ? next_data_22 : _GEN_85; // @[Regfile.scala 29:28 Regfile.scala 29:28]
  wire [31:0] _GEN_87 = 5'h17 == io_reg_read_1_op1_addr ? next_data_23 : _GEN_86; // @[Regfile.scala 29:28 Regfile.scala 29:28]
  wire [31:0] _GEN_88 = 5'h18 == io_reg_read_1_op1_addr ? next_data_24 : _GEN_87; // @[Regfile.scala 29:28 Regfile.scala 29:28]
  wire [31:0] _GEN_89 = 5'h19 == io_reg_read_1_op1_addr ? next_data_25 : _GEN_88; // @[Regfile.scala 29:28 Regfile.scala 29:28]
  wire [31:0] _GEN_90 = 5'h1a == io_reg_read_1_op1_addr ? next_data_26 : _GEN_89; // @[Regfile.scala 29:28 Regfile.scala 29:28]
  wire [31:0] _GEN_91 = 5'h1b == io_reg_read_1_op1_addr ? next_data_27 : _GEN_90; // @[Regfile.scala 29:28 Regfile.scala 29:28]
  wire [31:0] _GEN_92 = 5'h1c == io_reg_read_1_op1_addr ? next_data_28 : _GEN_91; // @[Regfile.scala 29:28 Regfile.scala 29:28]
  wire [31:0] _GEN_93 = 5'h1d == io_reg_read_1_op1_addr ? next_data_29 : _GEN_92; // @[Regfile.scala 29:28 Regfile.scala 29:28]
  wire [31:0] _GEN_94 = 5'h1e == io_reg_read_1_op1_addr ? next_data_30 : _GEN_93; // @[Regfile.scala 29:28 Regfile.scala 29:28]
  wire [31:0] _GEN_97 = 5'h1 == io_reg_read_1_op2_addr ? next_data_1 : 32'h0; // @[Regfile.scala 30:28 Regfile.scala 30:28]
  wire [31:0] _GEN_98 = 5'h2 == io_reg_read_1_op2_addr ? next_data_2 : _GEN_97; // @[Regfile.scala 30:28 Regfile.scala 30:28]
  wire [31:0] _GEN_99 = 5'h3 == io_reg_read_1_op2_addr ? next_data_3 : _GEN_98; // @[Regfile.scala 30:28 Regfile.scala 30:28]
  wire [31:0] _GEN_100 = 5'h4 == io_reg_read_1_op2_addr ? next_data_4 : _GEN_99; // @[Regfile.scala 30:28 Regfile.scala 30:28]
  wire [31:0] _GEN_101 = 5'h5 == io_reg_read_1_op2_addr ? next_data_5 : _GEN_100; // @[Regfile.scala 30:28 Regfile.scala 30:28]
  wire [31:0] _GEN_102 = 5'h6 == io_reg_read_1_op2_addr ? next_data_6 : _GEN_101; // @[Regfile.scala 30:28 Regfile.scala 30:28]
  wire [31:0] _GEN_103 = 5'h7 == io_reg_read_1_op2_addr ? next_data_7 : _GEN_102; // @[Regfile.scala 30:28 Regfile.scala 30:28]
  wire [31:0] _GEN_104 = 5'h8 == io_reg_read_1_op2_addr ? next_data_8 : _GEN_103; // @[Regfile.scala 30:28 Regfile.scala 30:28]
  wire [31:0] _GEN_105 = 5'h9 == io_reg_read_1_op2_addr ? next_data_9 : _GEN_104; // @[Regfile.scala 30:28 Regfile.scala 30:28]
  wire [31:0] _GEN_106 = 5'ha == io_reg_read_1_op2_addr ? next_data_10 : _GEN_105; // @[Regfile.scala 30:28 Regfile.scala 30:28]
  wire [31:0] _GEN_107 = 5'hb == io_reg_read_1_op2_addr ? next_data_11 : _GEN_106; // @[Regfile.scala 30:28 Regfile.scala 30:28]
  wire [31:0] _GEN_108 = 5'hc == io_reg_read_1_op2_addr ? next_data_12 : _GEN_107; // @[Regfile.scala 30:28 Regfile.scala 30:28]
  wire [31:0] _GEN_109 = 5'hd == io_reg_read_1_op2_addr ? next_data_13 : _GEN_108; // @[Regfile.scala 30:28 Regfile.scala 30:28]
  wire [31:0] _GEN_110 = 5'he == io_reg_read_1_op2_addr ? next_data_14 : _GEN_109; // @[Regfile.scala 30:28 Regfile.scala 30:28]
  wire [31:0] _GEN_111 = 5'hf == io_reg_read_1_op2_addr ? next_data_15 : _GEN_110; // @[Regfile.scala 30:28 Regfile.scala 30:28]
  wire [31:0] _GEN_112 = 5'h10 == io_reg_read_1_op2_addr ? next_data_16 : _GEN_111; // @[Regfile.scala 30:28 Regfile.scala 30:28]
  wire [31:0] _GEN_113 = 5'h11 == io_reg_read_1_op2_addr ? next_data_17 : _GEN_112; // @[Regfile.scala 30:28 Regfile.scala 30:28]
  wire [31:0] _GEN_114 = 5'h12 == io_reg_read_1_op2_addr ? next_data_18 : _GEN_113; // @[Regfile.scala 30:28 Regfile.scala 30:28]
  wire [31:0] _GEN_115 = 5'h13 == io_reg_read_1_op2_addr ? next_data_19 : _GEN_114; // @[Regfile.scala 30:28 Regfile.scala 30:28]
  wire [31:0] _GEN_116 = 5'h14 == io_reg_read_1_op2_addr ? next_data_20 : _GEN_115; // @[Regfile.scala 30:28 Regfile.scala 30:28]
  wire [31:0] _GEN_117 = 5'h15 == io_reg_read_1_op2_addr ? next_data_21 : _GEN_116; // @[Regfile.scala 30:28 Regfile.scala 30:28]
  wire [31:0] _GEN_118 = 5'h16 == io_reg_read_1_op2_addr ? next_data_22 : _GEN_117; // @[Regfile.scala 30:28 Regfile.scala 30:28]
  wire [31:0] _GEN_119 = 5'h17 == io_reg_read_1_op2_addr ? next_data_23 : _GEN_118; // @[Regfile.scala 30:28 Regfile.scala 30:28]
  wire [31:0] _GEN_120 = 5'h18 == io_reg_read_1_op2_addr ? next_data_24 : _GEN_119; // @[Regfile.scala 30:28 Regfile.scala 30:28]
  wire [31:0] _GEN_121 = 5'h19 == io_reg_read_1_op2_addr ? next_data_25 : _GEN_120; // @[Regfile.scala 30:28 Regfile.scala 30:28]
  wire [31:0] _GEN_122 = 5'h1a == io_reg_read_1_op2_addr ? next_data_26 : _GEN_121; // @[Regfile.scala 30:28 Regfile.scala 30:28]
  wire [31:0] _GEN_123 = 5'h1b == io_reg_read_1_op2_addr ? next_data_27 : _GEN_122; // @[Regfile.scala 30:28 Regfile.scala 30:28]
  wire [31:0] _GEN_124 = 5'h1c == io_reg_read_1_op2_addr ? next_data_28 : _GEN_123; // @[Regfile.scala 30:28 Regfile.scala 30:28]
  wire [31:0] _GEN_125 = 5'h1d == io_reg_read_1_op2_addr ? next_data_29 : _GEN_124; // @[Regfile.scala 30:28 Regfile.scala 30:28]
  wire [31:0] _GEN_126 = 5'h1e == io_reg_read_1_op2_addr ? next_data_30 : _GEN_125; // @[Regfile.scala 30:28 Regfile.scala 30:28]
  assign io_reg_read_0_op1_data = 5'h1f == io_reg_read_0_op1_addr ? next_data_31 : _GEN_30; // @[Regfile.scala 29:28 Regfile.scala 29:28]
  assign io_reg_read_0_op2_data = 5'h1f == io_reg_read_0_op2_addr ? next_data_31 : _GEN_62; // @[Regfile.scala 30:28 Regfile.scala 30:28]
  assign io_reg_read_1_op1_data = 5'h1f == io_reg_read_1_op1_addr ? next_data_31 : _GEN_94; // @[Regfile.scala 29:28 Regfile.scala 29:28]
  assign io_reg_read_1_op2_data = 5'h1f == io_reg_read_1_op2_addr ? next_data_31 : _GEN_126; // @[Regfile.scala 30:28 Regfile.scala 30:28]
  always @(posedge clock) begin
    if (reset) begin // @[Regfile.scala 18:24]
      regfile_1 <= 32'h0; // @[Regfile.scala 18:24]
    end else if (io_rob_commit_i_1_valid & commit_idx_1[1]) begin // @[Regfile.scala 25:93]
      regfile_1 <= io_rob_commit_i_1_bits_commit_data;
    end else if (io_rob_commit_i_0_valid & commit_idx_0[1]) begin // @[Regfile.scala 25:93]
      regfile_1 <= io_rob_commit_i_0_bits_commit_data;
    end
    if (reset) begin // @[Regfile.scala 18:24]
      regfile_2 <= 32'h0; // @[Regfile.scala 18:24]
    end else if (io_rob_commit_i_1_valid & commit_idx_1[2]) begin // @[Regfile.scala 25:93]
      regfile_2 <= io_rob_commit_i_1_bits_commit_data;
    end else if (io_rob_commit_i_0_valid & commit_idx_0[2]) begin // @[Regfile.scala 25:93]
      regfile_2 <= io_rob_commit_i_0_bits_commit_data;
    end
    if (reset) begin // @[Regfile.scala 18:24]
      regfile_3 <= 32'h0; // @[Regfile.scala 18:24]
    end else if (io_rob_commit_i_1_valid & commit_idx_1[3]) begin // @[Regfile.scala 25:93]
      regfile_3 <= io_rob_commit_i_1_bits_commit_data;
    end else if (io_rob_commit_i_0_valid & commit_idx_0[3]) begin // @[Regfile.scala 25:93]
      regfile_3 <= io_rob_commit_i_0_bits_commit_data;
    end
    if (reset) begin // @[Regfile.scala 18:24]
      regfile_4 <= 32'h0; // @[Regfile.scala 18:24]
    end else if (io_rob_commit_i_1_valid & commit_idx_1[4]) begin // @[Regfile.scala 25:93]
      regfile_4 <= io_rob_commit_i_1_bits_commit_data;
    end else if (io_rob_commit_i_0_valid & commit_idx_0[4]) begin // @[Regfile.scala 25:93]
      regfile_4 <= io_rob_commit_i_0_bits_commit_data;
    end
    if (reset) begin // @[Regfile.scala 18:24]
      regfile_5 <= 32'h0; // @[Regfile.scala 18:24]
    end else if (io_rob_commit_i_1_valid & commit_idx_1[5]) begin // @[Regfile.scala 25:93]
      regfile_5 <= io_rob_commit_i_1_bits_commit_data;
    end else if (io_rob_commit_i_0_valid & commit_idx_0[5]) begin // @[Regfile.scala 25:93]
      regfile_5 <= io_rob_commit_i_0_bits_commit_data;
    end
    if (reset) begin // @[Regfile.scala 18:24]
      regfile_6 <= 32'h0; // @[Regfile.scala 18:24]
    end else if (io_rob_commit_i_1_valid & commit_idx_1[6]) begin // @[Regfile.scala 25:93]
      regfile_6 <= io_rob_commit_i_1_bits_commit_data;
    end else if (io_rob_commit_i_0_valid & commit_idx_0[6]) begin // @[Regfile.scala 25:93]
      regfile_6 <= io_rob_commit_i_0_bits_commit_data;
    end
    if (reset) begin // @[Regfile.scala 18:24]
      regfile_7 <= 32'h0; // @[Regfile.scala 18:24]
    end else if (io_rob_commit_i_1_valid & commit_idx_1[7]) begin // @[Regfile.scala 25:93]
      regfile_7 <= io_rob_commit_i_1_bits_commit_data;
    end else if (io_rob_commit_i_0_valid & commit_idx_0[7]) begin // @[Regfile.scala 25:93]
      regfile_7 <= io_rob_commit_i_0_bits_commit_data;
    end
    if (reset) begin // @[Regfile.scala 18:24]
      regfile_8 <= 32'h0; // @[Regfile.scala 18:24]
    end else if (io_rob_commit_i_1_valid & commit_idx_1[8]) begin // @[Regfile.scala 25:93]
      regfile_8 <= io_rob_commit_i_1_bits_commit_data;
    end else if (io_rob_commit_i_0_valid & commit_idx_0[8]) begin // @[Regfile.scala 25:93]
      regfile_8 <= io_rob_commit_i_0_bits_commit_data;
    end
    if (reset) begin // @[Regfile.scala 18:24]
      regfile_9 <= 32'h0; // @[Regfile.scala 18:24]
    end else if (io_rob_commit_i_1_valid & commit_idx_1[9]) begin // @[Regfile.scala 25:93]
      regfile_9 <= io_rob_commit_i_1_bits_commit_data;
    end else if (io_rob_commit_i_0_valid & commit_idx_0[9]) begin // @[Regfile.scala 25:93]
      regfile_9 <= io_rob_commit_i_0_bits_commit_data;
    end
    if (reset) begin // @[Regfile.scala 18:24]
      regfile_10 <= 32'h0; // @[Regfile.scala 18:24]
    end else if (io_rob_commit_i_1_valid & commit_idx_1[10]) begin // @[Regfile.scala 25:93]
      regfile_10 <= io_rob_commit_i_1_bits_commit_data;
    end else if (io_rob_commit_i_0_valid & commit_idx_0[10]) begin // @[Regfile.scala 25:93]
      regfile_10 <= io_rob_commit_i_0_bits_commit_data;
    end
    if (reset) begin // @[Regfile.scala 18:24]
      regfile_11 <= 32'h0; // @[Regfile.scala 18:24]
    end else if (io_rob_commit_i_1_valid & commit_idx_1[11]) begin // @[Regfile.scala 25:93]
      regfile_11 <= io_rob_commit_i_1_bits_commit_data;
    end else if (io_rob_commit_i_0_valid & commit_idx_0[11]) begin // @[Regfile.scala 25:93]
      regfile_11 <= io_rob_commit_i_0_bits_commit_data;
    end
    if (reset) begin // @[Regfile.scala 18:24]
      regfile_12 <= 32'h0; // @[Regfile.scala 18:24]
    end else if (io_rob_commit_i_1_valid & commit_idx_1[12]) begin // @[Regfile.scala 25:93]
      regfile_12 <= io_rob_commit_i_1_bits_commit_data;
    end else if (io_rob_commit_i_0_valid & commit_idx_0[12]) begin // @[Regfile.scala 25:93]
      regfile_12 <= io_rob_commit_i_0_bits_commit_data;
    end
    if (reset) begin // @[Regfile.scala 18:24]
      regfile_13 <= 32'h0; // @[Regfile.scala 18:24]
    end else if (io_rob_commit_i_1_valid & commit_idx_1[13]) begin // @[Regfile.scala 25:93]
      regfile_13 <= io_rob_commit_i_1_bits_commit_data;
    end else if (io_rob_commit_i_0_valid & commit_idx_0[13]) begin // @[Regfile.scala 25:93]
      regfile_13 <= io_rob_commit_i_0_bits_commit_data;
    end
    if (reset) begin // @[Regfile.scala 18:24]
      regfile_14 <= 32'h0; // @[Regfile.scala 18:24]
    end else if (io_rob_commit_i_1_valid & commit_idx_1[14]) begin // @[Regfile.scala 25:93]
      regfile_14 <= io_rob_commit_i_1_bits_commit_data;
    end else if (io_rob_commit_i_0_valid & commit_idx_0[14]) begin // @[Regfile.scala 25:93]
      regfile_14 <= io_rob_commit_i_0_bits_commit_data;
    end
    if (reset) begin // @[Regfile.scala 18:24]
      regfile_15 <= 32'h0; // @[Regfile.scala 18:24]
    end else if (io_rob_commit_i_1_valid & commit_idx_1[15]) begin // @[Regfile.scala 25:93]
      regfile_15 <= io_rob_commit_i_1_bits_commit_data;
    end else if (io_rob_commit_i_0_valid & commit_idx_0[15]) begin // @[Regfile.scala 25:93]
      regfile_15 <= io_rob_commit_i_0_bits_commit_data;
    end
    if (reset) begin // @[Regfile.scala 18:24]
      regfile_16 <= 32'h0; // @[Regfile.scala 18:24]
    end else if (io_rob_commit_i_1_valid & commit_idx_1[16]) begin // @[Regfile.scala 25:93]
      regfile_16 <= io_rob_commit_i_1_bits_commit_data;
    end else if (io_rob_commit_i_0_valid & commit_idx_0[16]) begin // @[Regfile.scala 25:93]
      regfile_16 <= io_rob_commit_i_0_bits_commit_data;
    end
    if (reset) begin // @[Regfile.scala 18:24]
      regfile_17 <= 32'h0; // @[Regfile.scala 18:24]
    end else if (io_rob_commit_i_1_valid & commit_idx_1[17]) begin // @[Regfile.scala 25:93]
      regfile_17 <= io_rob_commit_i_1_bits_commit_data;
    end else if (io_rob_commit_i_0_valid & commit_idx_0[17]) begin // @[Regfile.scala 25:93]
      regfile_17 <= io_rob_commit_i_0_bits_commit_data;
    end
    if (reset) begin // @[Regfile.scala 18:24]
      regfile_18 <= 32'h0; // @[Regfile.scala 18:24]
    end else if (io_rob_commit_i_1_valid & commit_idx_1[18]) begin // @[Regfile.scala 25:93]
      regfile_18 <= io_rob_commit_i_1_bits_commit_data;
    end else if (io_rob_commit_i_0_valid & commit_idx_0[18]) begin // @[Regfile.scala 25:93]
      regfile_18 <= io_rob_commit_i_0_bits_commit_data;
    end
    if (reset) begin // @[Regfile.scala 18:24]
      regfile_19 <= 32'h0; // @[Regfile.scala 18:24]
    end else if (io_rob_commit_i_1_valid & commit_idx_1[19]) begin // @[Regfile.scala 25:93]
      regfile_19 <= io_rob_commit_i_1_bits_commit_data;
    end else if (io_rob_commit_i_0_valid & commit_idx_0[19]) begin // @[Regfile.scala 25:93]
      regfile_19 <= io_rob_commit_i_0_bits_commit_data;
    end
    if (reset) begin // @[Regfile.scala 18:24]
      regfile_20 <= 32'h0; // @[Regfile.scala 18:24]
    end else if (io_rob_commit_i_1_valid & commit_idx_1[20]) begin // @[Regfile.scala 25:93]
      regfile_20 <= io_rob_commit_i_1_bits_commit_data;
    end else if (io_rob_commit_i_0_valid & commit_idx_0[20]) begin // @[Regfile.scala 25:93]
      regfile_20 <= io_rob_commit_i_0_bits_commit_data;
    end
    if (reset) begin // @[Regfile.scala 18:24]
      regfile_21 <= 32'h0; // @[Regfile.scala 18:24]
    end else if (io_rob_commit_i_1_valid & commit_idx_1[21]) begin // @[Regfile.scala 25:93]
      regfile_21 <= io_rob_commit_i_1_bits_commit_data;
    end else if (io_rob_commit_i_0_valid & commit_idx_0[21]) begin // @[Regfile.scala 25:93]
      regfile_21 <= io_rob_commit_i_0_bits_commit_data;
    end
    if (reset) begin // @[Regfile.scala 18:24]
      regfile_22 <= 32'h0; // @[Regfile.scala 18:24]
    end else if (io_rob_commit_i_1_valid & commit_idx_1[22]) begin // @[Regfile.scala 25:93]
      regfile_22 <= io_rob_commit_i_1_bits_commit_data;
    end else if (io_rob_commit_i_0_valid & commit_idx_0[22]) begin // @[Regfile.scala 25:93]
      regfile_22 <= io_rob_commit_i_0_bits_commit_data;
    end
    if (reset) begin // @[Regfile.scala 18:24]
      regfile_23 <= 32'h0; // @[Regfile.scala 18:24]
    end else if (io_rob_commit_i_1_valid & commit_idx_1[23]) begin // @[Regfile.scala 25:93]
      regfile_23 <= io_rob_commit_i_1_bits_commit_data;
    end else if (io_rob_commit_i_0_valid & commit_idx_0[23]) begin // @[Regfile.scala 25:93]
      regfile_23 <= io_rob_commit_i_0_bits_commit_data;
    end
    if (reset) begin // @[Regfile.scala 18:24]
      regfile_24 <= 32'h0; // @[Regfile.scala 18:24]
    end else if (io_rob_commit_i_1_valid & commit_idx_1[24]) begin // @[Regfile.scala 25:93]
      regfile_24 <= io_rob_commit_i_1_bits_commit_data;
    end else if (io_rob_commit_i_0_valid & commit_idx_0[24]) begin // @[Regfile.scala 25:93]
      regfile_24 <= io_rob_commit_i_0_bits_commit_data;
    end
    if (reset) begin // @[Regfile.scala 18:24]
      regfile_25 <= 32'h0; // @[Regfile.scala 18:24]
    end else if (io_rob_commit_i_1_valid & commit_idx_1[25]) begin // @[Regfile.scala 25:93]
      regfile_25 <= io_rob_commit_i_1_bits_commit_data;
    end else if (io_rob_commit_i_0_valid & commit_idx_0[25]) begin // @[Regfile.scala 25:93]
      regfile_25 <= io_rob_commit_i_0_bits_commit_data;
    end
    if (reset) begin // @[Regfile.scala 18:24]
      regfile_26 <= 32'h0; // @[Regfile.scala 18:24]
    end else if (io_rob_commit_i_1_valid & commit_idx_1[26]) begin // @[Regfile.scala 25:93]
      regfile_26 <= io_rob_commit_i_1_bits_commit_data;
    end else if (io_rob_commit_i_0_valid & commit_idx_0[26]) begin // @[Regfile.scala 25:93]
      regfile_26 <= io_rob_commit_i_0_bits_commit_data;
    end
    if (reset) begin // @[Regfile.scala 18:24]
      regfile_27 <= 32'h0; // @[Regfile.scala 18:24]
    end else if (io_rob_commit_i_1_valid & commit_idx_1[27]) begin // @[Regfile.scala 25:93]
      regfile_27 <= io_rob_commit_i_1_bits_commit_data;
    end else if (io_rob_commit_i_0_valid & commit_idx_0[27]) begin // @[Regfile.scala 25:93]
      regfile_27 <= io_rob_commit_i_0_bits_commit_data;
    end
    if (reset) begin // @[Regfile.scala 18:24]
      regfile_28 <= 32'h0; // @[Regfile.scala 18:24]
    end else if (io_rob_commit_i_1_valid & commit_idx_1[28]) begin // @[Regfile.scala 25:93]
      regfile_28 <= io_rob_commit_i_1_bits_commit_data;
    end else if (io_rob_commit_i_0_valid & commit_idx_0[28]) begin // @[Regfile.scala 25:93]
      regfile_28 <= io_rob_commit_i_0_bits_commit_data;
    end
    if (reset) begin // @[Regfile.scala 18:24]
      regfile_29 <= 32'h0; // @[Regfile.scala 18:24]
    end else if (io_rob_commit_i_1_valid & commit_idx_1[29]) begin // @[Regfile.scala 25:93]
      regfile_29 <= io_rob_commit_i_1_bits_commit_data;
    end else if (io_rob_commit_i_0_valid & commit_idx_0[29]) begin // @[Regfile.scala 25:93]
      regfile_29 <= io_rob_commit_i_0_bits_commit_data;
    end
    if (reset) begin // @[Regfile.scala 18:24]
      regfile_30 <= 32'h0; // @[Regfile.scala 18:24]
    end else if (io_rob_commit_i_1_valid & commit_idx_1[30]) begin // @[Regfile.scala 25:93]
      regfile_30 <= io_rob_commit_i_1_bits_commit_data;
    end else if (io_rob_commit_i_0_valid & commit_idx_0[30]) begin // @[Regfile.scala 25:93]
      regfile_30 <= io_rob_commit_i_0_bits_commit_data;
    end
    if (reset) begin // @[Regfile.scala 18:24]
      regfile_31 <= 32'h0; // @[Regfile.scala 18:24]
    end else if (io_rob_commit_i_1_valid & commit_idx_1[31]) begin // @[Regfile.scala 25:93]
      regfile_31 <= io_rob_commit_i_1_bits_commit_data;
    end else if (io_rob_commit_i_0_valid & commit_idx_0[31]) begin // @[Regfile.scala 25:93]
      regfile_31 <= io_rob_commit_i_0_bits_commit_data;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  regfile_1 = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  regfile_2 = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  regfile_3 = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  regfile_4 = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  regfile_5 = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  regfile_6 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  regfile_7 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  regfile_8 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  regfile_9 = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  regfile_10 = _RAND_9[31:0];
  _RAND_10 = {1{`RANDOM}};
  regfile_11 = _RAND_10[31:0];
  _RAND_11 = {1{`RANDOM}};
  regfile_12 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  regfile_13 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  regfile_14 = _RAND_13[31:0];
  _RAND_14 = {1{`RANDOM}};
  regfile_15 = _RAND_14[31:0];
  _RAND_15 = {1{`RANDOM}};
  regfile_16 = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  regfile_17 = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  regfile_18 = _RAND_17[31:0];
  _RAND_18 = {1{`RANDOM}};
  regfile_19 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  regfile_20 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  regfile_21 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  regfile_22 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  regfile_23 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  regfile_24 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  regfile_25 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  regfile_26 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  regfile_27 = _RAND_26[31:0];
  _RAND_27 = {1{`RANDOM}};
  regfile_28 = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  regfile_29 = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  regfile_30 = _RAND_29[31:0];
  _RAND_30 = {1{`RANDOM}};
  regfile_31 = _RAND_30[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Rob(
  input         clock,
  input         reset,
  input         io_rob_allocate_allocate_req_valid,
  input         io_rob_allocate_allocate_req_bits_0,
  input         io_rob_allocate_allocate_req_bits_1,
  input         io_rob_allocate_allocate_info_valid,
  input  [2:0]  io_rob_allocate_allocate_info_bits_0_rob_idx,
  input         io_rob_allocate_allocate_info_bits_0_inst_valid,
  input  [31:0] io_rob_allocate_allocate_info_bits_0_inst_addr,
  input  [5:0]  io_rob_allocate_allocate_info_bits_0_uop,
  input  [2:0]  io_rob_allocate_allocate_info_bits_0_unit_sel,
  input         io_rob_allocate_allocate_info_bits_0_need_imm,
  input  [31:0] io_rob_allocate_allocate_info_bits_0_commit_addr,
  input  [3:0]  io_rob_allocate_allocate_info_bits_0_gh_info,
  input  [31:0] io_rob_allocate_allocate_info_bits_0_imm_data,
  input         io_rob_allocate_allocate_info_bits_0_flush_on_commit,
  input         io_rob_allocate_allocate_info_bits_0_predict_taken,
  input  [2:0]  io_rob_allocate_allocate_info_bits_1_rob_idx,
  input         io_rob_allocate_allocate_info_bits_1_inst_valid,
  input  [31:0] io_rob_allocate_allocate_info_bits_1_inst_addr,
  input  [5:0]  io_rob_allocate_allocate_info_bits_1_uop,
  input  [2:0]  io_rob_allocate_allocate_info_bits_1_unit_sel,
  input         io_rob_allocate_allocate_info_bits_1_need_imm,
  input  [31:0] io_rob_allocate_allocate_info_bits_1_commit_addr,
  input  [3:0]  io_rob_allocate_allocate_info_bits_1_gh_info,
  input  [31:0] io_rob_allocate_allocate_info_bits_1_imm_data,
  input         io_rob_allocate_allocate_info_bits_1_flush_on_commit,
  input         io_rob_allocate_allocate_info_bits_1_predict_taken,
  output        io_rob_allocate_allocate_resp_valid,
  output [2:0]  io_rob_allocate_allocate_resp_bits_rob_idx_0,
  output [2:0]  io_rob_allocate_allocate_resp_bits_rob_idx_1,
  output        io_rob_allocate_allocate_resp_bits_enq_valid_mask_0,
  output        io_rob_allocate_allocate_resp_bits_enq_valid_mask_1,
  input         io_rob_init_info_valid,
  input         io_rob_init_info_bits_0_is_valid,
  input  [2:0]  io_rob_init_info_bits_0_des_rob,
  input  [2:0]  io_rob_init_info_bits_0_op1_rob,
  input  [2:0]  io_rob_init_info_bits_0_op2_rob,
  input  [31:0] io_rob_init_info_bits_0_op1_regData,
  input  [31:0] io_rob_init_info_bits_0_op2_regData,
  input         io_rob_init_info_bits_0_op1_in_rob,
  input         io_rob_init_info_bits_0_op2_in_rob,
  input         io_rob_init_info_bits_1_is_valid,
  input  [2:0]  io_rob_init_info_bits_1_des_rob,
  input  [2:0]  io_rob_init_info_bits_1_op1_rob,
  input  [2:0]  io_rob_init_info_bits_1_op2_rob,
  input  [31:0] io_rob_init_info_bits_1_op1_regData,
  input  [31:0] io_rob_init_info_bits_1_op2_regData,
  input         io_rob_init_info_bits_1_op1_in_rob,
  input         io_rob_init_info_bits_1_op2_in_rob,
  input         io_wb_info_i_0_valid,
  input  [2:0]  io_wb_info_i_0_bits_rob_idx,
  input  [31:0] io_wb_info_i_0_bits_data,
  input         io_wb_info_i_1_valid,
  input  [2:0]  io_wb_info_i_1_bits_rob_idx,
  input  [31:0] io_wb_info_i_1_bits_data,
  input         io_wb_info_i_2_valid,
  input  [2:0]  io_wb_info_i_2_bits_rob_idx,
  input  [31:0] io_wb_info_i_2_bits_data,
  input  [31:0] io_wb_info_i_2_bits_target_addr,
  input         io_wb_info_i_2_bits_is_taken,
  input         io_wb_info_i_2_bits_predict_miss,
  input         io_wb_info_i_3_valid,
  input  [2:0]  io_wb_info_i_3_bits_rob_idx,
  input  [31:0] io_wb_info_i_3_bits_data,
  input         io_wb_info_i_4_valid,
  input  [2:0]  io_wb_info_i_4_bits_rob_idx,
  input  [31:0] io_wb_info_i_4_bits_data,
  output        io_dispatch_info_o_0_valid,
  output [5:0]  io_dispatch_info_o_0_bits_uop,
  output        io_dispatch_info_o_0_bits_need_imm,
  output [2:0]  io_dispatch_info_o_0_bits_rob_idx,
  output [31:0] io_dispatch_info_o_0_bits_op1_data,
  output [31:0] io_dispatch_info_o_0_bits_op2_data,
  output [31:0] io_dispatch_info_o_0_bits_imm_data,
  output        io_dispatch_info_o_1_valid,
  output [5:0]  io_dispatch_info_o_1_bits_uop,
  output        io_dispatch_info_o_1_bits_need_imm,
  output [2:0]  io_dispatch_info_o_1_bits_rob_idx,
  output [31:0] io_dispatch_info_o_1_bits_op1_data,
  output [31:0] io_dispatch_info_o_1_bits_op2_data,
  output [31:0] io_dispatch_info_o_1_bits_imm_data,
  output        io_dispatch_info_o_2_valid,
  output [5:0]  io_dispatch_info_o_2_bits_uop,
  output [2:0]  io_dispatch_info_o_2_bits_rob_idx,
  output [31:0] io_dispatch_info_o_2_bits_inst_addr,
  output [31:0] io_dispatch_info_o_2_bits_op1_data,
  output [31:0] io_dispatch_info_o_2_bits_op2_data,
  output [31:0] io_dispatch_info_o_2_bits_imm_data,
  output        io_dispatch_info_o_2_bits_predict_taken,
  output        io_dispatch_info_o_3_valid,
  output [2:0]  io_dispatch_info_o_3_bits_rob_idx,
  output [31:0] io_dispatch_info_o_3_bits_op1_data,
  output [31:0] io_dispatch_info_o_3_bits_op2_data,
  input         io_dispatch_info_o_4_ready,
  output        io_dispatch_info_o_4_valid,
  output [5:0]  io_dispatch_info_o_4_bits_uop,
  output [2:0]  io_dispatch_info_o_4_bits_rob_idx,
  output [31:0] io_dispatch_info_o_4_bits_op1_data,
  output [31:0] io_dispatch_info_o_4_bits_op2_data,
  output [31:0] io_dispatch_info_o_4_bits_imm_data,
  output        io_rob_commit_0_valid,
  output [2:0]  io_rob_commit_0_bits_des_rob,
  output [4:0]  io_rob_commit_0_bits_commit_addr,
  output [31:0] io_rob_commit_0_bits_commit_data,
  output        io_rob_commit_1_valid,
  output [2:0]  io_rob_commit_1_bits_des_rob,
  output [4:0]  io_rob_commit_1_bits_commit_addr,
  output [31:0] io_rob_commit_1_bits_commit_data,
  output        io_branch_info_valid,
  output [31:0] io_branch_info_bits_target_addr,
  output [31:0] io_branch_info_bits_inst_addr,
  output [3:0]  io_branch_info_bits_gh_update,
  output        io_branch_info_bits_is_branch,
  output        io_branch_info_bits_is_taken,
  output        io_branch_info_bits_predict_miss,
  output        io_need_flush
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [31:0] _RAND_86;
  reg [31:0] _RAND_87;
  reg [31:0] _RAND_88;
  reg [31:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [31:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
  reg [31:0] _RAND_118;
  reg [31:0] _RAND_119;
  reg [31:0] _RAND_120;
  reg [31:0] _RAND_121;
  reg [31:0] _RAND_122;
  reg [31:0] _RAND_123;
  reg [31:0] _RAND_124;
  reg [31:0] _RAND_125;
  reg [31:0] _RAND_126;
  reg [31:0] _RAND_127;
  reg [31:0] _RAND_128;
  reg [31:0] _RAND_129;
  reg [31:0] _RAND_130;
  reg [31:0] _RAND_131;
  reg [31:0] _RAND_132;
  reg [31:0] _RAND_133;
  reg [31:0] _RAND_134;
  reg [31:0] _RAND_135;
  reg [31:0] _RAND_136;
  reg [31:0] _RAND_137;
  reg [31:0] _RAND_138;
  reg [31:0] _RAND_139;
  reg [31:0] _RAND_140;
  reg [31:0] _RAND_141;
  reg [31:0] _RAND_142;
  reg [31:0] _RAND_143;
  reg [31:0] _RAND_144;
  reg [31:0] _RAND_145;
  reg [31:0] _RAND_146;
  reg [31:0] _RAND_147;
  reg [31:0] _RAND_148;
  reg [31:0] _RAND_149;
  reg [31:0] _RAND_150;
  reg [31:0] _RAND_151;
  reg [31:0] _RAND_152;
  reg [31:0] _RAND_153;
  reg [31:0] _RAND_154;
  reg [31:0] _RAND_155;
  reg [31:0] _RAND_156;
  reg [31:0] _RAND_157;
  reg [31:0] _RAND_158;
  reg [31:0] _RAND_159;
  reg [31:0] _RAND_160;
  reg [31:0] _RAND_161;
  reg [31:0] _RAND_162;
  reg [31:0] _RAND_163;
  reg [31:0] _RAND_164;
  reg [31:0] _RAND_165;
  reg [31:0] _RAND_166;
  reg [31:0] _RAND_167;
  reg [31:0] _RAND_168;
  reg [31:0] _RAND_169;
  reg [31:0] _RAND_170;
  reg [31:0] _RAND_171;
  reg [31:0] _RAND_172;
  reg [31:0] _RAND_173;
  reg [31:0] _RAND_174;
  reg [31:0] _RAND_175;
  reg [31:0] _RAND_176;
  reg [31:0] _RAND_177;
  reg [31:0] _RAND_178;
  reg [31:0] _RAND_179;
  reg [31:0] _RAND_180;
  reg [31:0] _RAND_181;
  reg [31:0] _RAND_182;
  reg [31:0] _RAND_183;
  reg [31:0] _RAND_184;
  reg [31:0] _RAND_185;
  reg [31:0] _RAND_186;
  reg [31:0] _RAND_187;
  reg [31:0] _RAND_188;
  reg [31:0] _RAND_189;
  reg [31:0] _RAND_190;
  reg [31:0] _RAND_191;
  reg [31:0] _RAND_192;
  reg [31:0] _RAND_193;
  reg [31:0] _RAND_194;
  reg [31:0] _RAND_195;
  reg [31:0] _RAND_196;
  reg [31:0] _RAND_197;
  reg [31:0] _RAND_198;
  reg [31:0] _RAND_199;
  reg [31:0] _RAND_200;
  reg [31:0] _RAND_201;
  reg [31:0] _RAND_202;
  reg [31:0] _RAND_203;
`endif // RANDOMIZE_REG_INIT
  reg  rob_info_0_is_valid; // @[Rob.scala 175:27]
  reg  rob_info_0_busy; // @[Rob.scala 175:27]
  reg [5:0] rob_info_0_uop; // @[Rob.scala 175:27]
  reg [2:0] rob_info_0_unit_sel; // @[Rob.scala 175:27]
  reg  rob_info_0_need_imm; // @[Rob.scala 175:27]
  reg [31:0] rob_info_0_inst_addr; // @[Rob.scala 175:27]
  reg [4:0] rob_info_0_commit_addr; // @[Rob.scala 175:27]
  reg [31:0] rob_info_0_commit_data; // @[Rob.scala 175:27]
  reg  rob_info_0_commit_ready; // @[Rob.scala 175:27]
  reg  rob_info_0_is_branch; // @[Rob.scala 175:27]
  reg  rob_info_0_predict_taken; // @[Rob.scala 175:27]
  reg  rob_info_0_is_taken; // @[Rob.scala 175:27]
  reg  rob_info_0_predict_miss; // @[Rob.scala 175:27]
  reg [3:0] rob_info_0_gh_info; // @[Rob.scala 175:27]
  reg  rob_info_0_op1_ready; // @[Rob.scala 175:27]
  reg [2:0] rob_info_0_op1_tag; // @[Rob.scala 175:27]
  reg [31:0] rob_info_0_op1_data; // @[Rob.scala 175:27]
  reg  rob_info_0_op2_ready; // @[Rob.scala 175:27]
  reg [2:0] rob_info_0_op2_tag; // @[Rob.scala 175:27]
  reg [31:0] rob_info_0_op2_data; // @[Rob.scala 175:27]
  reg [31:0] rob_info_0_imm_data; // @[Rob.scala 175:27]
  reg  rob_info_0_is_init; // @[Rob.scala 175:27]
  reg  rob_info_0_flush_on_commit; // @[Rob.scala 175:27]
  reg  rob_info_1_is_valid; // @[Rob.scala 175:27]
  reg  rob_info_1_busy; // @[Rob.scala 175:27]
  reg [5:0] rob_info_1_uop; // @[Rob.scala 175:27]
  reg [2:0] rob_info_1_unit_sel; // @[Rob.scala 175:27]
  reg  rob_info_1_need_imm; // @[Rob.scala 175:27]
  reg [31:0] rob_info_1_inst_addr; // @[Rob.scala 175:27]
  reg [4:0] rob_info_1_commit_addr; // @[Rob.scala 175:27]
  reg [31:0] rob_info_1_commit_data; // @[Rob.scala 175:27]
  reg  rob_info_1_commit_ready; // @[Rob.scala 175:27]
  reg  rob_info_1_is_branch; // @[Rob.scala 175:27]
  reg  rob_info_1_predict_taken; // @[Rob.scala 175:27]
  reg  rob_info_1_is_taken; // @[Rob.scala 175:27]
  reg  rob_info_1_predict_miss; // @[Rob.scala 175:27]
  reg [3:0] rob_info_1_gh_info; // @[Rob.scala 175:27]
  reg  rob_info_1_op1_ready; // @[Rob.scala 175:27]
  reg [2:0] rob_info_1_op1_tag; // @[Rob.scala 175:27]
  reg [31:0] rob_info_1_op1_data; // @[Rob.scala 175:27]
  reg  rob_info_1_op2_ready; // @[Rob.scala 175:27]
  reg [2:0] rob_info_1_op2_tag; // @[Rob.scala 175:27]
  reg [31:0] rob_info_1_op2_data; // @[Rob.scala 175:27]
  reg [31:0] rob_info_1_imm_data; // @[Rob.scala 175:27]
  reg  rob_info_1_is_init; // @[Rob.scala 175:27]
  reg  rob_info_1_flush_on_commit; // @[Rob.scala 175:27]
  reg  rob_info_2_is_valid; // @[Rob.scala 175:27]
  reg  rob_info_2_busy; // @[Rob.scala 175:27]
  reg [5:0] rob_info_2_uop; // @[Rob.scala 175:27]
  reg [2:0] rob_info_2_unit_sel; // @[Rob.scala 175:27]
  reg  rob_info_2_need_imm; // @[Rob.scala 175:27]
  reg [31:0] rob_info_2_inst_addr; // @[Rob.scala 175:27]
  reg [4:0] rob_info_2_commit_addr; // @[Rob.scala 175:27]
  reg [31:0] rob_info_2_commit_data; // @[Rob.scala 175:27]
  reg  rob_info_2_commit_ready; // @[Rob.scala 175:27]
  reg  rob_info_2_is_branch; // @[Rob.scala 175:27]
  reg  rob_info_2_predict_taken; // @[Rob.scala 175:27]
  reg  rob_info_2_is_taken; // @[Rob.scala 175:27]
  reg  rob_info_2_predict_miss; // @[Rob.scala 175:27]
  reg [3:0] rob_info_2_gh_info; // @[Rob.scala 175:27]
  reg  rob_info_2_op1_ready; // @[Rob.scala 175:27]
  reg [2:0] rob_info_2_op1_tag; // @[Rob.scala 175:27]
  reg [31:0] rob_info_2_op1_data; // @[Rob.scala 175:27]
  reg  rob_info_2_op2_ready; // @[Rob.scala 175:27]
  reg [2:0] rob_info_2_op2_tag; // @[Rob.scala 175:27]
  reg [31:0] rob_info_2_op2_data; // @[Rob.scala 175:27]
  reg [31:0] rob_info_2_imm_data; // @[Rob.scala 175:27]
  reg  rob_info_2_is_init; // @[Rob.scala 175:27]
  reg  rob_info_2_flush_on_commit; // @[Rob.scala 175:27]
  reg  rob_info_3_is_valid; // @[Rob.scala 175:27]
  reg  rob_info_3_busy; // @[Rob.scala 175:27]
  reg [5:0] rob_info_3_uop; // @[Rob.scala 175:27]
  reg [2:0] rob_info_3_unit_sel; // @[Rob.scala 175:27]
  reg  rob_info_3_need_imm; // @[Rob.scala 175:27]
  reg [31:0] rob_info_3_inst_addr; // @[Rob.scala 175:27]
  reg [4:0] rob_info_3_commit_addr; // @[Rob.scala 175:27]
  reg [31:0] rob_info_3_commit_data; // @[Rob.scala 175:27]
  reg  rob_info_3_commit_ready; // @[Rob.scala 175:27]
  reg  rob_info_3_is_branch; // @[Rob.scala 175:27]
  reg  rob_info_3_predict_taken; // @[Rob.scala 175:27]
  reg  rob_info_3_is_taken; // @[Rob.scala 175:27]
  reg  rob_info_3_predict_miss; // @[Rob.scala 175:27]
  reg [3:0] rob_info_3_gh_info; // @[Rob.scala 175:27]
  reg  rob_info_3_op1_ready; // @[Rob.scala 175:27]
  reg [2:0] rob_info_3_op1_tag; // @[Rob.scala 175:27]
  reg [31:0] rob_info_3_op1_data; // @[Rob.scala 175:27]
  reg  rob_info_3_op2_ready; // @[Rob.scala 175:27]
  reg [2:0] rob_info_3_op2_tag; // @[Rob.scala 175:27]
  reg [31:0] rob_info_3_op2_data; // @[Rob.scala 175:27]
  reg [31:0] rob_info_3_imm_data; // @[Rob.scala 175:27]
  reg  rob_info_3_is_init; // @[Rob.scala 175:27]
  reg  rob_info_3_flush_on_commit; // @[Rob.scala 175:27]
  reg  rob_info_4_is_valid; // @[Rob.scala 175:27]
  reg  rob_info_4_busy; // @[Rob.scala 175:27]
  reg [5:0] rob_info_4_uop; // @[Rob.scala 175:27]
  reg [2:0] rob_info_4_unit_sel; // @[Rob.scala 175:27]
  reg  rob_info_4_need_imm; // @[Rob.scala 175:27]
  reg [31:0] rob_info_4_inst_addr; // @[Rob.scala 175:27]
  reg [4:0] rob_info_4_commit_addr; // @[Rob.scala 175:27]
  reg [31:0] rob_info_4_commit_data; // @[Rob.scala 175:27]
  reg  rob_info_4_commit_ready; // @[Rob.scala 175:27]
  reg  rob_info_4_is_branch; // @[Rob.scala 175:27]
  reg  rob_info_4_predict_taken; // @[Rob.scala 175:27]
  reg  rob_info_4_is_taken; // @[Rob.scala 175:27]
  reg  rob_info_4_predict_miss; // @[Rob.scala 175:27]
  reg [3:0] rob_info_4_gh_info; // @[Rob.scala 175:27]
  reg  rob_info_4_op1_ready; // @[Rob.scala 175:27]
  reg [2:0] rob_info_4_op1_tag; // @[Rob.scala 175:27]
  reg [31:0] rob_info_4_op1_data; // @[Rob.scala 175:27]
  reg  rob_info_4_op2_ready; // @[Rob.scala 175:27]
  reg [2:0] rob_info_4_op2_tag; // @[Rob.scala 175:27]
  reg [31:0] rob_info_4_op2_data; // @[Rob.scala 175:27]
  reg [31:0] rob_info_4_imm_data; // @[Rob.scala 175:27]
  reg  rob_info_4_is_init; // @[Rob.scala 175:27]
  reg  rob_info_4_flush_on_commit; // @[Rob.scala 175:27]
  reg  rob_info_5_is_valid; // @[Rob.scala 175:27]
  reg  rob_info_5_busy; // @[Rob.scala 175:27]
  reg [5:0] rob_info_5_uop; // @[Rob.scala 175:27]
  reg [2:0] rob_info_5_unit_sel; // @[Rob.scala 175:27]
  reg  rob_info_5_need_imm; // @[Rob.scala 175:27]
  reg [31:0] rob_info_5_inst_addr; // @[Rob.scala 175:27]
  reg [4:0] rob_info_5_commit_addr; // @[Rob.scala 175:27]
  reg [31:0] rob_info_5_commit_data; // @[Rob.scala 175:27]
  reg  rob_info_5_commit_ready; // @[Rob.scala 175:27]
  reg  rob_info_5_is_branch; // @[Rob.scala 175:27]
  reg  rob_info_5_predict_taken; // @[Rob.scala 175:27]
  reg  rob_info_5_is_taken; // @[Rob.scala 175:27]
  reg  rob_info_5_predict_miss; // @[Rob.scala 175:27]
  reg [3:0] rob_info_5_gh_info; // @[Rob.scala 175:27]
  reg  rob_info_5_op1_ready; // @[Rob.scala 175:27]
  reg [2:0] rob_info_5_op1_tag; // @[Rob.scala 175:27]
  reg [31:0] rob_info_5_op1_data; // @[Rob.scala 175:27]
  reg  rob_info_5_op2_ready; // @[Rob.scala 175:27]
  reg [2:0] rob_info_5_op2_tag; // @[Rob.scala 175:27]
  reg [31:0] rob_info_5_op2_data; // @[Rob.scala 175:27]
  reg [31:0] rob_info_5_imm_data; // @[Rob.scala 175:27]
  reg  rob_info_5_is_init; // @[Rob.scala 175:27]
  reg  rob_info_5_flush_on_commit; // @[Rob.scala 175:27]
  reg  rob_info_6_is_valid; // @[Rob.scala 175:27]
  reg  rob_info_6_busy; // @[Rob.scala 175:27]
  reg [5:0] rob_info_6_uop; // @[Rob.scala 175:27]
  reg [2:0] rob_info_6_unit_sel; // @[Rob.scala 175:27]
  reg  rob_info_6_need_imm; // @[Rob.scala 175:27]
  reg [31:0] rob_info_6_inst_addr; // @[Rob.scala 175:27]
  reg [4:0] rob_info_6_commit_addr; // @[Rob.scala 175:27]
  reg [31:0] rob_info_6_commit_data; // @[Rob.scala 175:27]
  reg  rob_info_6_commit_ready; // @[Rob.scala 175:27]
  reg  rob_info_6_is_branch; // @[Rob.scala 175:27]
  reg  rob_info_6_predict_taken; // @[Rob.scala 175:27]
  reg  rob_info_6_is_taken; // @[Rob.scala 175:27]
  reg  rob_info_6_predict_miss; // @[Rob.scala 175:27]
  reg [3:0] rob_info_6_gh_info; // @[Rob.scala 175:27]
  reg  rob_info_6_op1_ready; // @[Rob.scala 175:27]
  reg [2:0] rob_info_6_op1_tag; // @[Rob.scala 175:27]
  reg [31:0] rob_info_6_op1_data; // @[Rob.scala 175:27]
  reg  rob_info_6_op2_ready; // @[Rob.scala 175:27]
  reg [2:0] rob_info_6_op2_tag; // @[Rob.scala 175:27]
  reg [31:0] rob_info_6_op2_data; // @[Rob.scala 175:27]
  reg [31:0] rob_info_6_imm_data; // @[Rob.scala 175:27]
  reg  rob_info_6_is_init; // @[Rob.scala 175:27]
  reg  rob_info_6_flush_on_commit; // @[Rob.scala 175:27]
  reg  rob_info_7_is_valid; // @[Rob.scala 175:27]
  reg  rob_info_7_busy; // @[Rob.scala 175:27]
  reg [5:0] rob_info_7_uop; // @[Rob.scala 175:27]
  reg [2:0] rob_info_7_unit_sel; // @[Rob.scala 175:27]
  reg  rob_info_7_need_imm; // @[Rob.scala 175:27]
  reg [31:0] rob_info_7_inst_addr; // @[Rob.scala 175:27]
  reg [4:0] rob_info_7_commit_addr; // @[Rob.scala 175:27]
  reg [31:0] rob_info_7_commit_data; // @[Rob.scala 175:27]
  reg  rob_info_7_commit_ready; // @[Rob.scala 175:27]
  reg  rob_info_7_is_branch; // @[Rob.scala 175:27]
  reg  rob_info_7_predict_taken; // @[Rob.scala 175:27]
  reg  rob_info_7_is_taken; // @[Rob.scala 175:27]
  reg  rob_info_7_predict_miss; // @[Rob.scala 175:27]
  reg [3:0] rob_info_7_gh_info; // @[Rob.scala 175:27]
  reg  rob_info_7_op1_ready; // @[Rob.scala 175:27]
  reg [2:0] rob_info_7_op1_tag; // @[Rob.scala 175:27]
  reg [31:0] rob_info_7_op1_data; // @[Rob.scala 175:27]
  reg  rob_info_7_op2_ready; // @[Rob.scala 175:27]
  reg [2:0] rob_info_7_op2_tag; // @[Rob.scala 175:27]
  reg [31:0] rob_info_7_op2_data; // @[Rob.scala 175:27]
  reg [31:0] rob_info_7_imm_data; // @[Rob.scala 175:27]
  reg  rob_info_7_is_init; // @[Rob.scala 175:27]
  reg  rob_info_7_flush_on_commit; // @[Rob.scala 175:27]
  reg [7:0] head; // @[Rob.scala 176:31]
  reg [7:0] tail; // @[Rob.scala 178:31]
  reg  maybe_full; // @[Rob.scala 179:31]
  wire  hit_head = head == tail; // @[Rob.scala 180:29]
  wire  is_empty = hit_head & ~maybe_full; // @[Rob.scala 182:33]
  wire  might_hit_head_mask_0 = tail == head & ~is_empty; // @[Rob.scala 193:48]
  wire  inst_valid_mask_0 = io_rob_allocate_allocate_req_bits_0 & io_rob_allocate_allocate_req_valid; // @[Rob.scala 186:64]
  wire  _T_4 = ~might_hit_head_mask_0; // @[Rob.scala 195:42]
  wire [6:0] hi = tail[6:0]; // @[Rob.scala 167:12]
  wire  lo = tail[7]; // @[Rob.scala 167:29]
  wire [7:0] _T_6 = {hi,lo}; // @[Cat.scala 30:58]
  wire [7:0] enq_idxs_1 = inst_valid_mask_0 & ~might_hit_head_mask_0 ? _T_6 : tail; // @[Rob.scala 195:20]
  wire  might_hit_1 = might_hit_head_mask_0 | enq_idxs_1 == head & ~is_empty; // @[Rob.scala 193:27]
  wire  inst_valid_mask_1 = io_rob_allocate_allocate_req_bits_1 & io_rob_allocate_allocate_req_valid; // @[Rob.scala 186:64]
  reg  waiting_delay; // @[Rob.scala 187:30]
  reg  need_flush; // @[Rob.scala 188:27]
  wire  _T_11 = ~might_hit_1; // @[Rob.scala 195:42]
  wire [6:0] hi_1 = enq_idxs_1[6:0]; // @[Rob.scala 167:12]
  wire  lo_1 = enq_idxs_1[7]; // @[Rob.scala 167:29]
  wire [7:0] _T_13 = {hi_1,lo_1}; // @[Cat.scala 30:58]
  wire  enq_valid_mask_0 = _T_4 & inst_valid_mask_0; // @[Rob.scala 197:79]
  wire  enq_valid_mask_1 = _T_11 & inst_valid_mask_1; // @[Rob.scala 197:79]
  wire  do_enq = enq_valid_mask_0 | enq_valid_mask_1; // @[Rob.scala 198:43]
  wire [3:0] hi_2 = tail[7:4]; // @[OneHot.scala 30:18]
  wire [3:0] lo_2 = tail[3:0]; // @[OneHot.scala 31:18]
  wire  hi_3 = |hi_2; // @[OneHot.scala 32:14]
  wire [3:0] _T_14 = hi_2 | lo_2; // @[OneHot.scala 32:28]
  wire [1:0] hi_4 = _T_14[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] lo_3 = _T_14[1:0]; // @[OneHot.scala 31:18]
  wire  hi_5 = |hi_4; // @[OneHot.scala 32:14]
  wire [1:0] _T_15 = hi_4 | lo_3; // @[OneHot.scala 32:28]
  wire  lo_4 = _T_15[1]; // @[CircuitMath.scala 30:8]
  wire [1:0] lo_5 = {hi_5,lo_4}; // @[Cat.scala 30:58]
  wire [3:0] hi_6 = enq_idxs_1[7:4]; // @[OneHot.scala 30:18]
  wire [3:0] lo_6 = enq_idxs_1[3:0]; // @[OneHot.scala 31:18]
  wire  hi_7 = |hi_6; // @[OneHot.scala 32:14]
  wire [3:0] _T_17 = hi_6 | lo_6; // @[OneHot.scala 32:28]
  wire [1:0] hi_8 = _T_17[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] lo_7 = _T_17[1:0]; // @[OneHot.scala 31:18]
  wire  hi_9 = |hi_8; // @[OneHot.scala 32:14]
  wire [1:0] _T_18 = hi_8 | lo_7; // @[OneHot.scala 32:28]
  wire  lo_8 = _T_18[1]; // @[CircuitMath.scala 30:8]
  wire [1:0] lo_9 = {hi_9,lo_8}; // @[Cat.scala 30:58]
  wire [3:0] dispatch_idxs_hi = head[7:4]; // @[OneHot.scala 30:18]
  wire [3:0] dispatch_idxs_lo = head[3:0]; // @[OneHot.scala 31:18]
  wire  dispatch_idxs_hi_1 = |dispatch_idxs_hi; // @[OneHot.scala 32:14]
  wire [3:0] _dispatch_idxs_T = dispatch_idxs_hi | dispatch_idxs_lo; // @[OneHot.scala 32:28]
  wire [1:0] dispatch_idxs_hi_2 = _dispatch_idxs_T[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] dispatch_idxs_lo_1 = _dispatch_idxs_T[1:0]; // @[OneHot.scala 31:18]
  wire  dispatch_idxs_hi_3 = |dispatch_idxs_hi_2; // @[OneHot.scala 32:14]
  wire [1:0] _dispatch_idxs_T_1 = dispatch_idxs_hi_2 | dispatch_idxs_lo_1; // @[OneHot.scala 32:28]
  wire  dispatch_idxs_lo_2 = _dispatch_idxs_T_1[1]; // @[CircuitMath.scala 30:8]
  wire [2:0] dispatch_idxs_0 = {dispatch_idxs_hi_1,dispatch_idxs_hi_3,dispatch_idxs_lo_2}; // @[Cat.scala 30:58]
  wire [6:0] dispatch_idxs_hi_4 = head[6:0]; // @[Rob.scala 167:12]
  wire  dispatch_idxs_lo_4 = head[7]; // @[Rob.scala 167:29]
  wire [7:0] _dispatch_idxs_T_3 = {dispatch_idxs_hi_4,dispatch_idxs_lo_4}; // @[Cat.scala 30:58]
  wire [3:0] dispatch_idxs_hi_5 = _dispatch_idxs_T_3[7:4]; // @[OneHot.scala 30:18]
  wire [3:0] dispatch_idxs_lo_5 = _dispatch_idxs_T_3[3:0]; // @[OneHot.scala 31:18]
  wire  dispatch_idxs_hi_6 = |dispatch_idxs_hi_5; // @[OneHot.scala 32:14]
  wire [3:0] _dispatch_idxs_T_4 = dispatch_idxs_hi_5 | dispatch_idxs_lo_5; // @[OneHot.scala 32:28]
  wire [1:0] dispatch_idxs_hi_7 = _dispatch_idxs_T_4[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] dispatch_idxs_lo_6 = _dispatch_idxs_T_4[1:0]; // @[OneHot.scala 31:18]
  wire  dispatch_idxs_hi_8 = |dispatch_idxs_hi_7; // @[OneHot.scala 32:14]
  wire [1:0] _dispatch_idxs_T_5 = dispatch_idxs_hi_7 | dispatch_idxs_lo_6; // @[OneHot.scala 32:28]
  wire  dispatch_idxs_lo_7 = _dispatch_idxs_T_5[1]; // @[CircuitMath.scala 30:8]
  wire [2:0] dispatch_idxs_1 = {dispatch_idxs_hi_6,dispatch_idxs_hi_8,dispatch_idxs_lo_7}; // @[Cat.scala 30:58]
  wire [5:0] dispatch_idxs_hi_9 = head[5:0]; // @[Rob.scala 167:12]
  wire [1:0] dispatch_idxs_lo_9 = head[7:6]; // @[Rob.scala 167:29]
  wire [7:0] _dispatch_idxs_T_7 = {dispatch_idxs_hi_9,dispatch_idxs_lo_9}; // @[Cat.scala 30:58]
  wire [3:0] dispatch_idxs_hi_10 = _dispatch_idxs_T_7[7:4]; // @[OneHot.scala 30:18]
  wire [3:0] dispatch_idxs_lo_10 = _dispatch_idxs_T_7[3:0]; // @[OneHot.scala 31:18]
  wire  dispatch_idxs_hi_11 = |dispatch_idxs_hi_10; // @[OneHot.scala 32:14]
  wire [3:0] _dispatch_idxs_T_8 = dispatch_idxs_hi_10 | dispatch_idxs_lo_10; // @[OneHot.scala 32:28]
  wire [1:0] dispatch_idxs_hi_12 = _dispatch_idxs_T_8[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] dispatch_idxs_lo_11 = _dispatch_idxs_T_8[1:0]; // @[OneHot.scala 31:18]
  wire  dispatch_idxs_hi_13 = |dispatch_idxs_hi_12; // @[OneHot.scala 32:14]
  wire [1:0] _dispatch_idxs_T_9 = dispatch_idxs_hi_12 | dispatch_idxs_lo_11; // @[OneHot.scala 32:28]
  wire  dispatch_idxs_lo_12 = _dispatch_idxs_T_9[1]; // @[CircuitMath.scala 30:8]
  wire [2:0] dispatch_idxs_2 = {dispatch_idxs_hi_11,dispatch_idxs_hi_13,dispatch_idxs_lo_12}; // @[Cat.scala 30:58]
  wire [4:0] dispatch_idxs_hi_14 = head[4:0]; // @[Rob.scala 167:12]
  wire [2:0] dispatch_idxs_lo_14 = head[7:5]; // @[Rob.scala 167:29]
  wire [7:0] _dispatch_idxs_T_11 = {dispatch_idxs_hi_14,dispatch_idxs_lo_14}; // @[Cat.scala 30:58]
  wire [3:0] dispatch_idxs_hi_15 = _dispatch_idxs_T_11[7:4]; // @[OneHot.scala 30:18]
  wire [3:0] dispatch_idxs_lo_15 = _dispatch_idxs_T_11[3:0]; // @[OneHot.scala 31:18]
  wire  dispatch_idxs_hi_16 = |dispatch_idxs_hi_15; // @[OneHot.scala 32:14]
  wire [3:0] _dispatch_idxs_T_12 = dispatch_idxs_hi_15 | dispatch_idxs_lo_15; // @[OneHot.scala 32:28]
  wire [1:0] dispatch_idxs_hi_17 = _dispatch_idxs_T_12[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] dispatch_idxs_lo_16 = _dispatch_idxs_T_12[1:0]; // @[OneHot.scala 31:18]
  wire  dispatch_idxs_hi_18 = |dispatch_idxs_hi_17; // @[OneHot.scala 32:14]
  wire [1:0] _dispatch_idxs_T_13 = dispatch_idxs_hi_17 | dispatch_idxs_lo_16; // @[OneHot.scala 32:28]
  wire  dispatch_idxs_lo_17 = _dispatch_idxs_T_13[1]; // @[CircuitMath.scala 30:8]
  wire [2:0] dispatch_idxs_3 = {dispatch_idxs_hi_16,dispatch_idxs_hi_18,dispatch_idxs_lo_17}; // @[Cat.scala 30:58]
  wire [7:0] _dispatch_idxs_T_15 = {dispatch_idxs_lo,dispatch_idxs_hi}; // @[Cat.scala 30:58]
  wire [3:0] dispatch_idxs_hi_20 = _dispatch_idxs_T_15[7:4]; // @[OneHot.scala 30:18]
  wire [3:0] dispatch_idxs_lo_20 = _dispatch_idxs_T_15[3:0]; // @[OneHot.scala 31:18]
  wire  dispatch_idxs_hi_21 = |dispatch_idxs_hi_20; // @[OneHot.scala 32:14]
  wire [3:0] _dispatch_idxs_T_16 = dispatch_idxs_hi_20 | dispatch_idxs_lo_20; // @[OneHot.scala 32:28]
  wire [1:0] dispatch_idxs_hi_22 = _dispatch_idxs_T_16[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] dispatch_idxs_lo_21 = _dispatch_idxs_T_16[1:0]; // @[OneHot.scala 31:18]
  wire  dispatch_idxs_hi_23 = |dispatch_idxs_hi_22; // @[OneHot.scala 32:14]
  wire [1:0] _dispatch_idxs_T_17 = dispatch_idxs_hi_22 | dispatch_idxs_lo_21; // @[OneHot.scala 32:28]
  wire  dispatch_idxs_lo_22 = _dispatch_idxs_T_17[1]; // @[CircuitMath.scala 30:8]
  wire [2:0] dispatch_idxs_4 = {dispatch_idxs_hi_21,dispatch_idxs_hi_23,dispatch_idxs_lo_22}; // @[Cat.scala 30:58]
  wire [2:0] dispatch_idxs_hi_24 = head[2:0]; // @[Rob.scala 167:12]
  wire [4:0] dispatch_idxs_lo_24 = head[7:3]; // @[Rob.scala 167:29]
  wire [7:0] _dispatch_idxs_T_19 = {dispatch_idxs_hi_24,dispatch_idxs_lo_24}; // @[Cat.scala 30:58]
  wire [3:0] dispatch_idxs_hi_25 = _dispatch_idxs_T_19[7:4]; // @[OneHot.scala 30:18]
  wire [3:0] dispatch_idxs_lo_25 = _dispatch_idxs_T_19[3:0]; // @[OneHot.scala 31:18]
  wire  dispatch_idxs_hi_26 = |dispatch_idxs_hi_25; // @[OneHot.scala 32:14]
  wire [3:0] _dispatch_idxs_T_20 = dispatch_idxs_hi_25 | dispatch_idxs_lo_25; // @[OneHot.scala 32:28]
  wire [1:0] dispatch_idxs_hi_27 = _dispatch_idxs_T_20[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] dispatch_idxs_lo_26 = _dispatch_idxs_T_20[1:0]; // @[OneHot.scala 31:18]
  wire  dispatch_idxs_hi_28 = |dispatch_idxs_hi_27; // @[OneHot.scala 32:14]
  wire [1:0] _dispatch_idxs_T_21 = dispatch_idxs_hi_27 | dispatch_idxs_lo_26; // @[OneHot.scala 32:28]
  wire  dispatch_idxs_lo_27 = _dispatch_idxs_T_21[1]; // @[CircuitMath.scala 30:8]
  wire [2:0] dispatch_idxs_5 = {dispatch_idxs_hi_26,dispatch_idxs_hi_28,dispatch_idxs_lo_27}; // @[Cat.scala 30:58]
  wire [1:0] dispatch_idxs_hi_29 = head[1:0]; // @[Rob.scala 167:12]
  wire [5:0] dispatch_idxs_lo_29 = head[7:2]; // @[Rob.scala 167:29]
  wire [7:0] _dispatch_idxs_T_23 = {dispatch_idxs_hi_29,dispatch_idxs_lo_29}; // @[Cat.scala 30:58]
  wire [3:0] dispatch_idxs_hi_30 = _dispatch_idxs_T_23[7:4]; // @[OneHot.scala 30:18]
  wire [3:0] dispatch_idxs_lo_30 = _dispatch_idxs_T_23[3:0]; // @[OneHot.scala 31:18]
  wire  dispatch_idxs_hi_31 = |dispatch_idxs_hi_30; // @[OneHot.scala 32:14]
  wire [3:0] _dispatch_idxs_T_24 = dispatch_idxs_hi_30 | dispatch_idxs_lo_30; // @[OneHot.scala 32:28]
  wire [1:0] dispatch_idxs_hi_32 = _dispatch_idxs_T_24[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] dispatch_idxs_lo_31 = _dispatch_idxs_T_24[1:0]; // @[OneHot.scala 31:18]
  wire  dispatch_idxs_hi_33 = |dispatch_idxs_hi_32; // @[OneHot.scala 32:14]
  wire [1:0] _dispatch_idxs_T_25 = dispatch_idxs_hi_32 | dispatch_idxs_lo_31; // @[OneHot.scala 32:28]
  wire  dispatch_idxs_lo_32 = _dispatch_idxs_T_25[1]; // @[CircuitMath.scala 30:8]
  wire [2:0] dispatch_idxs_6 = {dispatch_idxs_hi_31,dispatch_idxs_hi_33,dispatch_idxs_lo_32}; // @[Cat.scala 30:58]
  wire  dispatch_idxs_hi_34 = head[0]; // @[Rob.scala 167:12]
  wire [6:0] dispatch_idxs_lo_34 = head[7:1]; // @[Rob.scala 167:29]
  wire [7:0] _dispatch_idxs_T_27 = {dispatch_idxs_hi_34,dispatch_idxs_lo_34}; // @[Cat.scala 30:58]
  wire [3:0] dispatch_idxs_hi_35 = _dispatch_idxs_T_27[7:4]; // @[OneHot.scala 30:18]
  wire [3:0] dispatch_idxs_lo_35 = _dispatch_idxs_T_27[3:0]; // @[OneHot.scala 31:18]
  wire  dispatch_idxs_hi_36 = |dispatch_idxs_hi_35; // @[OneHot.scala 32:14]
  wire [3:0] _dispatch_idxs_T_28 = dispatch_idxs_hi_35 | dispatch_idxs_lo_35; // @[OneHot.scala 32:28]
  wire [1:0] dispatch_idxs_hi_37 = _dispatch_idxs_T_28[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] dispatch_idxs_lo_36 = _dispatch_idxs_T_28[1:0]; // @[OneHot.scala 31:18]
  wire  dispatch_idxs_hi_38 = |dispatch_idxs_hi_37; // @[OneHot.scala 32:14]
  wire [1:0] _dispatch_idxs_T_29 = dispatch_idxs_hi_37 | dispatch_idxs_lo_36; // @[OneHot.scala 32:28]
  wire  dispatch_idxs_lo_37 = _dispatch_idxs_T_29[1]; // @[CircuitMath.scala 30:8]
  wire [2:0] dispatch_idxs_7 = {dispatch_idxs_hi_36,dispatch_idxs_hi_38,dispatch_idxs_lo_37}; // @[Cat.scala 30:58]
  wire  _GEN_1 = 3'h1 == dispatch_idxs_0 ? rob_info_1_commit_ready : rob_info_0_commit_ready; // @[Rob.scala 211:54 Rob.scala 211:54]
  wire  _GEN_2 = 3'h2 == dispatch_idxs_0 ? rob_info_2_commit_ready : _GEN_1; // @[Rob.scala 211:54 Rob.scala 211:54]
  wire  _GEN_3 = 3'h3 == dispatch_idxs_0 ? rob_info_3_commit_ready : _GEN_2; // @[Rob.scala 211:54 Rob.scala 211:54]
  wire  _GEN_4 = 3'h4 == dispatch_idxs_0 ? rob_info_4_commit_ready : _GEN_3; // @[Rob.scala 211:54 Rob.scala 211:54]
  wire  _GEN_5 = 3'h5 == dispatch_idxs_0 ? rob_info_5_commit_ready : _GEN_4; // @[Rob.scala 211:54 Rob.scala 211:54]
  wire  _GEN_6 = 3'h6 == dispatch_idxs_0 ? rob_info_6_commit_ready : _GEN_5; // @[Rob.scala 211:54 Rob.scala 211:54]
  wire  _GEN_7 = 3'h7 == dispatch_idxs_0 ? rob_info_7_commit_ready : _GEN_6; // @[Rob.scala 211:54 Rob.scala 211:54]
  wire  _ready_mask_T = ~_GEN_7; // @[Rob.scala 211:54]
  wire  _GEN_9 = 3'h1 == dispatch_idxs_0 ? rob_info_1_busy : rob_info_0_busy; // @[Rob.scala 211:83 Rob.scala 211:83]
  wire  _GEN_10 = 3'h2 == dispatch_idxs_0 ? rob_info_2_busy : _GEN_9; // @[Rob.scala 211:83 Rob.scala 211:83]
  wire  _GEN_11 = 3'h3 == dispatch_idxs_0 ? rob_info_3_busy : _GEN_10; // @[Rob.scala 211:83 Rob.scala 211:83]
  wire  _GEN_12 = 3'h4 == dispatch_idxs_0 ? rob_info_4_busy : _GEN_11; // @[Rob.scala 211:83 Rob.scala 211:83]
  wire  _GEN_13 = 3'h5 == dispatch_idxs_0 ? rob_info_5_busy : _GEN_12; // @[Rob.scala 211:83 Rob.scala 211:83]
  wire  _GEN_14 = 3'h6 == dispatch_idxs_0 ? rob_info_6_busy : _GEN_13; // @[Rob.scala 211:83 Rob.scala 211:83]
  wire  _GEN_15 = 3'h7 == dispatch_idxs_0 ? rob_info_7_busy : _GEN_14; // @[Rob.scala 211:83 Rob.scala 211:83]
  wire  _ready_mask_T_1 = ~_GEN_15; // @[Rob.scala 211:83]
  wire  _GEN_17 = 3'h1 == dispatch_idxs_0 ? rob_info_1_is_valid : rob_info_0_is_valid; // @[Rob.scala 211:101 Rob.scala 211:101]
  wire  _GEN_18 = 3'h2 == dispatch_idxs_0 ? rob_info_2_is_valid : _GEN_17; // @[Rob.scala 211:101 Rob.scala 211:101]
  wire  _GEN_19 = 3'h3 == dispatch_idxs_0 ? rob_info_3_is_valid : _GEN_18; // @[Rob.scala 211:101 Rob.scala 211:101]
  wire  _GEN_20 = 3'h4 == dispatch_idxs_0 ? rob_info_4_is_valid : _GEN_19; // @[Rob.scala 211:101 Rob.scala 211:101]
  wire  _GEN_21 = 3'h5 == dispatch_idxs_0 ? rob_info_5_is_valid : _GEN_20; // @[Rob.scala 211:101 Rob.scala 211:101]
  wire  _GEN_22 = 3'h6 == dispatch_idxs_0 ? rob_info_6_is_valid : _GEN_21; // @[Rob.scala 211:101 Rob.scala 211:101]
  wire  _GEN_23 = 3'h7 == dispatch_idxs_0 ? rob_info_7_is_valid : _GEN_22; // @[Rob.scala 211:101 Rob.scala 211:101]
  wire  _GEN_25 = 3'h1 == dispatch_idxs_0 ? rob_info_1_op1_ready : rob_info_0_op1_ready; // @[Rob.scala 211:125 Rob.scala 211:125]
  wire  _GEN_26 = 3'h2 == dispatch_idxs_0 ? rob_info_2_op1_ready : _GEN_25; // @[Rob.scala 211:125 Rob.scala 211:125]
  wire  _GEN_27 = 3'h3 == dispatch_idxs_0 ? rob_info_3_op1_ready : _GEN_26; // @[Rob.scala 211:125 Rob.scala 211:125]
  wire  _GEN_28 = 3'h4 == dispatch_idxs_0 ? rob_info_4_op1_ready : _GEN_27; // @[Rob.scala 211:125 Rob.scala 211:125]
  wire  _GEN_29 = 3'h5 == dispatch_idxs_0 ? rob_info_5_op1_ready : _GEN_28; // @[Rob.scala 211:125 Rob.scala 211:125]
  wire  _GEN_30 = 3'h6 == dispatch_idxs_0 ? rob_info_6_op1_ready : _GEN_29; // @[Rob.scala 211:125 Rob.scala 211:125]
  wire  _GEN_31 = 3'h7 == dispatch_idxs_0 ? rob_info_7_op1_ready : _GEN_30; // @[Rob.scala 211:125 Rob.scala 211:125]
  wire  _GEN_33 = 3'h1 == dispatch_idxs_0 ? rob_info_1_op2_ready : rob_info_0_op2_ready; // @[Rob.scala 211:150 Rob.scala 211:150]
  wire  _GEN_34 = 3'h2 == dispatch_idxs_0 ? rob_info_2_op2_ready : _GEN_33; // @[Rob.scala 211:150 Rob.scala 211:150]
  wire  _GEN_35 = 3'h3 == dispatch_idxs_0 ? rob_info_3_op2_ready : _GEN_34; // @[Rob.scala 211:150 Rob.scala 211:150]
  wire  _GEN_36 = 3'h4 == dispatch_idxs_0 ? rob_info_4_op2_ready : _GEN_35; // @[Rob.scala 211:150 Rob.scala 211:150]
  wire  _GEN_37 = 3'h5 == dispatch_idxs_0 ? rob_info_5_op2_ready : _GEN_36; // @[Rob.scala 211:150 Rob.scala 211:150]
  wire  _GEN_38 = 3'h6 == dispatch_idxs_0 ? rob_info_6_op2_ready : _GEN_37; // @[Rob.scala 211:150 Rob.scala 211:150]
  wire  _GEN_39 = 3'h7 == dispatch_idxs_0 ? rob_info_7_op2_ready : _GEN_38; // @[Rob.scala 211:150 Rob.scala 211:150]
  wire  ready_mask_0 = ~_GEN_7 & ~_GEN_15 & _GEN_23 & _GEN_31 & _GEN_39; // @[Rob.scala 211:150]
  wire  _GEN_41 = 3'h1 == dispatch_idxs_1 ? rob_info_1_commit_ready : rob_info_0_commit_ready; // @[Rob.scala 211:54 Rob.scala 211:54]
  wire  _GEN_42 = 3'h2 == dispatch_idxs_1 ? rob_info_2_commit_ready : _GEN_41; // @[Rob.scala 211:54 Rob.scala 211:54]
  wire  _GEN_43 = 3'h3 == dispatch_idxs_1 ? rob_info_3_commit_ready : _GEN_42; // @[Rob.scala 211:54 Rob.scala 211:54]
  wire  _GEN_44 = 3'h4 == dispatch_idxs_1 ? rob_info_4_commit_ready : _GEN_43; // @[Rob.scala 211:54 Rob.scala 211:54]
  wire  _GEN_45 = 3'h5 == dispatch_idxs_1 ? rob_info_5_commit_ready : _GEN_44; // @[Rob.scala 211:54 Rob.scala 211:54]
  wire  _GEN_46 = 3'h6 == dispatch_idxs_1 ? rob_info_6_commit_ready : _GEN_45; // @[Rob.scala 211:54 Rob.scala 211:54]
  wire  _GEN_47 = 3'h7 == dispatch_idxs_1 ? rob_info_7_commit_ready : _GEN_46; // @[Rob.scala 211:54 Rob.scala 211:54]
  wire  _ready_mask_T_6 = ~_GEN_47; // @[Rob.scala 211:54]
  wire  _GEN_49 = 3'h1 == dispatch_idxs_1 ? rob_info_1_busy : rob_info_0_busy; // @[Rob.scala 211:83 Rob.scala 211:83]
  wire  _GEN_50 = 3'h2 == dispatch_idxs_1 ? rob_info_2_busy : _GEN_49; // @[Rob.scala 211:83 Rob.scala 211:83]
  wire  _GEN_51 = 3'h3 == dispatch_idxs_1 ? rob_info_3_busy : _GEN_50; // @[Rob.scala 211:83 Rob.scala 211:83]
  wire  _GEN_52 = 3'h4 == dispatch_idxs_1 ? rob_info_4_busy : _GEN_51; // @[Rob.scala 211:83 Rob.scala 211:83]
  wire  _GEN_53 = 3'h5 == dispatch_idxs_1 ? rob_info_5_busy : _GEN_52; // @[Rob.scala 211:83 Rob.scala 211:83]
  wire  _GEN_54 = 3'h6 == dispatch_idxs_1 ? rob_info_6_busy : _GEN_53; // @[Rob.scala 211:83 Rob.scala 211:83]
  wire  _GEN_55 = 3'h7 == dispatch_idxs_1 ? rob_info_7_busy : _GEN_54; // @[Rob.scala 211:83 Rob.scala 211:83]
  wire  _ready_mask_T_7 = ~_GEN_55; // @[Rob.scala 211:83]
  wire  _GEN_57 = 3'h1 == dispatch_idxs_1 ? rob_info_1_is_valid : rob_info_0_is_valid; // @[Rob.scala 211:101 Rob.scala 211:101]
  wire  _GEN_58 = 3'h2 == dispatch_idxs_1 ? rob_info_2_is_valid : _GEN_57; // @[Rob.scala 211:101 Rob.scala 211:101]
  wire  _GEN_59 = 3'h3 == dispatch_idxs_1 ? rob_info_3_is_valid : _GEN_58; // @[Rob.scala 211:101 Rob.scala 211:101]
  wire  _GEN_60 = 3'h4 == dispatch_idxs_1 ? rob_info_4_is_valid : _GEN_59; // @[Rob.scala 211:101 Rob.scala 211:101]
  wire  _GEN_61 = 3'h5 == dispatch_idxs_1 ? rob_info_5_is_valid : _GEN_60; // @[Rob.scala 211:101 Rob.scala 211:101]
  wire  _GEN_62 = 3'h6 == dispatch_idxs_1 ? rob_info_6_is_valid : _GEN_61; // @[Rob.scala 211:101 Rob.scala 211:101]
  wire  _GEN_63 = 3'h7 == dispatch_idxs_1 ? rob_info_7_is_valid : _GEN_62; // @[Rob.scala 211:101 Rob.scala 211:101]
  wire  _GEN_65 = 3'h1 == dispatch_idxs_1 ? rob_info_1_op1_ready : rob_info_0_op1_ready; // @[Rob.scala 211:125 Rob.scala 211:125]
  wire  _GEN_66 = 3'h2 == dispatch_idxs_1 ? rob_info_2_op1_ready : _GEN_65; // @[Rob.scala 211:125 Rob.scala 211:125]
  wire  _GEN_67 = 3'h3 == dispatch_idxs_1 ? rob_info_3_op1_ready : _GEN_66; // @[Rob.scala 211:125 Rob.scala 211:125]
  wire  _GEN_68 = 3'h4 == dispatch_idxs_1 ? rob_info_4_op1_ready : _GEN_67; // @[Rob.scala 211:125 Rob.scala 211:125]
  wire  _GEN_69 = 3'h5 == dispatch_idxs_1 ? rob_info_5_op1_ready : _GEN_68; // @[Rob.scala 211:125 Rob.scala 211:125]
  wire  _GEN_70 = 3'h6 == dispatch_idxs_1 ? rob_info_6_op1_ready : _GEN_69; // @[Rob.scala 211:125 Rob.scala 211:125]
  wire  _GEN_71 = 3'h7 == dispatch_idxs_1 ? rob_info_7_op1_ready : _GEN_70; // @[Rob.scala 211:125 Rob.scala 211:125]
  wire  _GEN_73 = 3'h1 == dispatch_idxs_1 ? rob_info_1_op2_ready : rob_info_0_op2_ready; // @[Rob.scala 211:150 Rob.scala 211:150]
  wire  _GEN_74 = 3'h2 == dispatch_idxs_1 ? rob_info_2_op2_ready : _GEN_73; // @[Rob.scala 211:150 Rob.scala 211:150]
  wire  _GEN_75 = 3'h3 == dispatch_idxs_1 ? rob_info_3_op2_ready : _GEN_74; // @[Rob.scala 211:150 Rob.scala 211:150]
  wire  _GEN_76 = 3'h4 == dispatch_idxs_1 ? rob_info_4_op2_ready : _GEN_75; // @[Rob.scala 211:150 Rob.scala 211:150]
  wire  _GEN_77 = 3'h5 == dispatch_idxs_1 ? rob_info_5_op2_ready : _GEN_76; // @[Rob.scala 211:150 Rob.scala 211:150]
  wire  _GEN_78 = 3'h6 == dispatch_idxs_1 ? rob_info_6_op2_ready : _GEN_77; // @[Rob.scala 211:150 Rob.scala 211:150]
  wire  _GEN_79 = 3'h7 == dispatch_idxs_1 ? rob_info_7_op2_ready : _GEN_78; // @[Rob.scala 211:150 Rob.scala 211:150]
  wire  ready_mask_1 = ~_GEN_47 & ~_GEN_55 & _GEN_63 & _GEN_71 & _GEN_79; // @[Rob.scala 211:150]
  wire  _GEN_81 = 3'h1 == dispatch_idxs_2 ? rob_info_1_commit_ready : rob_info_0_commit_ready; // @[Rob.scala 211:54 Rob.scala 211:54]
  wire  _GEN_82 = 3'h2 == dispatch_idxs_2 ? rob_info_2_commit_ready : _GEN_81; // @[Rob.scala 211:54 Rob.scala 211:54]
  wire  _GEN_83 = 3'h3 == dispatch_idxs_2 ? rob_info_3_commit_ready : _GEN_82; // @[Rob.scala 211:54 Rob.scala 211:54]
  wire  _GEN_84 = 3'h4 == dispatch_idxs_2 ? rob_info_4_commit_ready : _GEN_83; // @[Rob.scala 211:54 Rob.scala 211:54]
  wire  _GEN_85 = 3'h5 == dispatch_idxs_2 ? rob_info_5_commit_ready : _GEN_84; // @[Rob.scala 211:54 Rob.scala 211:54]
  wire  _GEN_86 = 3'h6 == dispatch_idxs_2 ? rob_info_6_commit_ready : _GEN_85; // @[Rob.scala 211:54 Rob.scala 211:54]
  wire  _GEN_87 = 3'h7 == dispatch_idxs_2 ? rob_info_7_commit_ready : _GEN_86; // @[Rob.scala 211:54 Rob.scala 211:54]
  wire  _ready_mask_T_12 = ~_GEN_87; // @[Rob.scala 211:54]
  wire  _GEN_89 = 3'h1 == dispatch_idxs_2 ? rob_info_1_busy : rob_info_0_busy; // @[Rob.scala 211:83 Rob.scala 211:83]
  wire  _GEN_90 = 3'h2 == dispatch_idxs_2 ? rob_info_2_busy : _GEN_89; // @[Rob.scala 211:83 Rob.scala 211:83]
  wire  _GEN_91 = 3'h3 == dispatch_idxs_2 ? rob_info_3_busy : _GEN_90; // @[Rob.scala 211:83 Rob.scala 211:83]
  wire  _GEN_92 = 3'h4 == dispatch_idxs_2 ? rob_info_4_busy : _GEN_91; // @[Rob.scala 211:83 Rob.scala 211:83]
  wire  _GEN_93 = 3'h5 == dispatch_idxs_2 ? rob_info_5_busy : _GEN_92; // @[Rob.scala 211:83 Rob.scala 211:83]
  wire  _GEN_94 = 3'h6 == dispatch_idxs_2 ? rob_info_6_busy : _GEN_93; // @[Rob.scala 211:83 Rob.scala 211:83]
  wire  _GEN_95 = 3'h7 == dispatch_idxs_2 ? rob_info_7_busy : _GEN_94; // @[Rob.scala 211:83 Rob.scala 211:83]
  wire  _ready_mask_T_13 = ~_GEN_95; // @[Rob.scala 211:83]
  wire  _GEN_97 = 3'h1 == dispatch_idxs_2 ? rob_info_1_is_valid : rob_info_0_is_valid; // @[Rob.scala 211:101 Rob.scala 211:101]
  wire  _GEN_98 = 3'h2 == dispatch_idxs_2 ? rob_info_2_is_valid : _GEN_97; // @[Rob.scala 211:101 Rob.scala 211:101]
  wire  _GEN_99 = 3'h3 == dispatch_idxs_2 ? rob_info_3_is_valid : _GEN_98; // @[Rob.scala 211:101 Rob.scala 211:101]
  wire  _GEN_100 = 3'h4 == dispatch_idxs_2 ? rob_info_4_is_valid : _GEN_99; // @[Rob.scala 211:101 Rob.scala 211:101]
  wire  _GEN_101 = 3'h5 == dispatch_idxs_2 ? rob_info_5_is_valid : _GEN_100; // @[Rob.scala 211:101 Rob.scala 211:101]
  wire  _GEN_102 = 3'h6 == dispatch_idxs_2 ? rob_info_6_is_valid : _GEN_101; // @[Rob.scala 211:101 Rob.scala 211:101]
  wire  _GEN_103 = 3'h7 == dispatch_idxs_2 ? rob_info_7_is_valid : _GEN_102; // @[Rob.scala 211:101 Rob.scala 211:101]
  wire  _GEN_105 = 3'h1 == dispatch_idxs_2 ? rob_info_1_op1_ready : rob_info_0_op1_ready; // @[Rob.scala 211:125 Rob.scala 211:125]
  wire  _GEN_106 = 3'h2 == dispatch_idxs_2 ? rob_info_2_op1_ready : _GEN_105; // @[Rob.scala 211:125 Rob.scala 211:125]
  wire  _GEN_107 = 3'h3 == dispatch_idxs_2 ? rob_info_3_op1_ready : _GEN_106; // @[Rob.scala 211:125 Rob.scala 211:125]
  wire  _GEN_108 = 3'h4 == dispatch_idxs_2 ? rob_info_4_op1_ready : _GEN_107; // @[Rob.scala 211:125 Rob.scala 211:125]
  wire  _GEN_109 = 3'h5 == dispatch_idxs_2 ? rob_info_5_op1_ready : _GEN_108; // @[Rob.scala 211:125 Rob.scala 211:125]
  wire  _GEN_110 = 3'h6 == dispatch_idxs_2 ? rob_info_6_op1_ready : _GEN_109; // @[Rob.scala 211:125 Rob.scala 211:125]
  wire  _GEN_111 = 3'h7 == dispatch_idxs_2 ? rob_info_7_op1_ready : _GEN_110; // @[Rob.scala 211:125 Rob.scala 211:125]
  wire  _GEN_113 = 3'h1 == dispatch_idxs_2 ? rob_info_1_op2_ready : rob_info_0_op2_ready; // @[Rob.scala 211:150 Rob.scala 211:150]
  wire  _GEN_114 = 3'h2 == dispatch_idxs_2 ? rob_info_2_op2_ready : _GEN_113; // @[Rob.scala 211:150 Rob.scala 211:150]
  wire  _GEN_115 = 3'h3 == dispatch_idxs_2 ? rob_info_3_op2_ready : _GEN_114; // @[Rob.scala 211:150 Rob.scala 211:150]
  wire  _GEN_116 = 3'h4 == dispatch_idxs_2 ? rob_info_4_op2_ready : _GEN_115; // @[Rob.scala 211:150 Rob.scala 211:150]
  wire  _GEN_117 = 3'h5 == dispatch_idxs_2 ? rob_info_5_op2_ready : _GEN_116; // @[Rob.scala 211:150 Rob.scala 211:150]
  wire  _GEN_118 = 3'h6 == dispatch_idxs_2 ? rob_info_6_op2_ready : _GEN_117; // @[Rob.scala 211:150 Rob.scala 211:150]
  wire  _GEN_119 = 3'h7 == dispatch_idxs_2 ? rob_info_7_op2_ready : _GEN_118; // @[Rob.scala 211:150 Rob.scala 211:150]
  wire  ready_mask_2 = ~_GEN_87 & ~_GEN_95 & _GEN_103 & _GEN_111 & _GEN_119; // @[Rob.scala 211:150]
  wire  _GEN_121 = 3'h1 == dispatch_idxs_3 ? rob_info_1_commit_ready : rob_info_0_commit_ready; // @[Rob.scala 211:54 Rob.scala 211:54]
  wire  _GEN_122 = 3'h2 == dispatch_idxs_3 ? rob_info_2_commit_ready : _GEN_121; // @[Rob.scala 211:54 Rob.scala 211:54]
  wire  _GEN_123 = 3'h3 == dispatch_idxs_3 ? rob_info_3_commit_ready : _GEN_122; // @[Rob.scala 211:54 Rob.scala 211:54]
  wire  _GEN_124 = 3'h4 == dispatch_idxs_3 ? rob_info_4_commit_ready : _GEN_123; // @[Rob.scala 211:54 Rob.scala 211:54]
  wire  _GEN_125 = 3'h5 == dispatch_idxs_3 ? rob_info_5_commit_ready : _GEN_124; // @[Rob.scala 211:54 Rob.scala 211:54]
  wire  _GEN_126 = 3'h6 == dispatch_idxs_3 ? rob_info_6_commit_ready : _GEN_125; // @[Rob.scala 211:54 Rob.scala 211:54]
  wire  _GEN_127 = 3'h7 == dispatch_idxs_3 ? rob_info_7_commit_ready : _GEN_126; // @[Rob.scala 211:54 Rob.scala 211:54]
  wire  _ready_mask_T_18 = ~_GEN_127; // @[Rob.scala 211:54]
  wire  _GEN_129 = 3'h1 == dispatch_idxs_3 ? rob_info_1_busy : rob_info_0_busy; // @[Rob.scala 211:83 Rob.scala 211:83]
  wire  _GEN_130 = 3'h2 == dispatch_idxs_3 ? rob_info_2_busy : _GEN_129; // @[Rob.scala 211:83 Rob.scala 211:83]
  wire  _GEN_131 = 3'h3 == dispatch_idxs_3 ? rob_info_3_busy : _GEN_130; // @[Rob.scala 211:83 Rob.scala 211:83]
  wire  _GEN_132 = 3'h4 == dispatch_idxs_3 ? rob_info_4_busy : _GEN_131; // @[Rob.scala 211:83 Rob.scala 211:83]
  wire  _GEN_133 = 3'h5 == dispatch_idxs_3 ? rob_info_5_busy : _GEN_132; // @[Rob.scala 211:83 Rob.scala 211:83]
  wire  _GEN_134 = 3'h6 == dispatch_idxs_3 ? rob_info_6_busy : _GEN_133; // @[Rob.scala 211:83 Rob.scala 211:83]
  wire  _GEN_135 = 3'h7 == dispatch_idxs_3 ? rob_info_7_busy : _GEN_134; // @[Rob.scala 211:83 Rob.scala 211:83]
  wire  _ready_mask_T_19 = ~_GEN_135; // @[Rob.scala 211:83]
  wire  _GEN_137 = 3'h1 == dispatch_idxs_3 ? rob_info_1_is_valid : rob_info_0_is_valid; // @[Rob.scala 211:101 Rob.scala 211:101]
  wire  _GEN_138 = 3'h2 == dispatch_idxs_3 ? rob_info_2_is_valid : _GEN_137; // @[Rob.scala 211:101 Rob.scala 211:101]
  wire  _GEN_139 = 3'h3 == dispatch_idxs_3 ? rob_info_3_is_valid : _GEN_138; // @[Rob.scala 211:101 Rob.scala 211:101]
  wire  _GEN_140 = 3'h4 == dispatch_idxs_3 ? rob_info_4_is_valid : _GEN_139; // @[Rob.scala 211:101 Rob.scala 211:101]
  wire  _GEN_141 = 3'h5 == dispatch_idxs_3 ? rob_info_5_is_valid : _GEN_140; // @[Rob.scala 211:101 Rob.scala 211:101]
  wire  _GEN_142 = 3'h6 == dispatch_idxs_3 ? rob_info_6_is_valid : _GEN_141; // @[Rob.scala 211:101 Rob.scala 211:101]
  wire  _GEN_143 = 3'h7 == dispatch_idxs_3 ? rob_info_7_is_valid : _GEN_142; // @[Rob.scala 211:101 Rob.scala 211:101]
  wire  _GEN_145 = 3'h1 == dispatch_idxs_3 ? rob_info_1_op1_ready : rob_info_0_op1_ready; // @[Rob.scala 211:125 Rob.scala 211:125]
  wire  _GEN_146 = 3'h2 == dispatch_idxs_3 ? rob_info_2_op1_ready : _GEN_145; // @[Rob.scala 211:125 Rob.scala 211:125]
  wire  _GEN_147 = 3'h3 == dispatch_idxs_3 ? rob_info_3_op1_ready : _GEN_146; // @[Rob.scala 211:125 Rob.scala 211:125]
  wire  _GEN_148 = 3'h4 == dispatch_idxs_3 ? rob_info_4_op1_ready : _GEN_147; // @[Rob.scala 211:125 Rob.scala 211:125]
  wire  _GEN_149 = 3'h5 == dispatch_idxs_3 ? rob_info_5_op1_ready : _GEN_148; // @[Rob.scala 211:125 Rob.scala 211:125]
  wire  _GEN_150 = 3'h6 == dispatch_idxs_3 ? rob_info_6_op1_ready : _GEN_149; // @[Rob.scala 211:125 Rob.scala 211:125]
  wire  _GEN_151 = 3'h7 == dispatch_idxs_3 ? rob_info_7_op1_ready : _GEN_150; // @[Rob.scala 211:125 Rob.scala 211:125]
  wire  _GEN_153 = 3'h1 == dispatch_idxs_3 ? rob_info_1_op2_ready : rob_info_0_op2_ready; // @[Rob.scala 211:150 Rob.scala 211:150]
  wire  _GEN_154 = 3'h2 == dispatch_idxs_3 ? rob_info_2_op2_ready : _GEN_153; // @[Rob.scala 211:150 Rob.scala 211:150]
  wire  _GEN_155 = 3'h3 == dispatch_idxs_3 ? rob_info_3_op2_ready : _GEN_154; // @[Rob.scala 211:150 Rob.scala 211:150]
  wire  _GEN_156 = 3'h4 == dispatch_idxs_3 ? rob_info_4_op2_ready : _GEN_155; // @[Rob.scala 211:150 Rob.scala 211:150]
  wire  _GEN_157 = 3'h5 == dispatch_idxs_3 ? rob_info_5_op2_ready : _GEN_156; // @[Rob.scala 211:150 Rob.scala 211:150]
  wire  _GEN_158 = 3'h6 == dispatch_idxs_3 ? rob_info_6_op2_ready : _GEN_157; // @[Rob.scala 211:150 Rob.scala 211:150]
  wire  _GEN_159 = 3'h7 == dispatch_idxs_3 ? rob_info_7_op2_ready : _GEN_158; // @[Rob.scala 211:150 Rob.scala 211:150]
  wire  ready_mask_3 = ~_GEN_127 & ~_GEN_135 & _GEN_143 & _GEN_151 & _GEN_159; // @[Rob.scala 211:150]
  wire  _GEN_161 = 3'h1 == dispatch_idxs_4 ? rob_info_1_commit_ready : rob_info_0_commit_ready; // @[Rob.scala 211:54 Rob.scala 211:54]
  wire  _GEN_162 = 3'h2 == dispatch_idxs_4 ? rob_info_2_commit_ready : _GEN_161; // @[Rob.scala 211:54 Rob.scala 211:54]
  wire  _GEN_163 = 3'h3 == dispatch_idxs_4 ? rob_info_3_commit_ready : _GEN_162; // @[Rob.scala 211:54 Rob.scala 211:54]
  wire  _GEN_164 = 3'h4 == dispatch_idxs_4 ? rob_info_4_commit_ready : _GEN_163; // @[Rob.scala 211:54 Rob.scala 211:54]
  wire  _GEN_165 = 3'h5 == dispatch_idxs_4 ? rob_info_5_commit_ready : _GEN_164; // @[Rob.scala 211:54 Rob.scala 211:54]
  wire  _GEN_166 = 3'h6 == dispatch_idxs_4 ? rob_info_6_commit_ready : _GEN_165; // @[Rob.scala 211:54 Rob.scala 211:54]
  wire  _GEN_167 = 3'h7 == dispatch_idxs_4 ? rob_info_7_commit_ready : _GEN_166; // @[Rob.scala 211:54 Rob.scala 211:54]
  wire  _ready_mask_T_24 = ~_GEN_167; // @[Rob.scala 211:54]
  wire  _GEN_169 = 3'h1 == dispatch_idxs_4 ? rob_info_1_busy : rob_info_0_busy; // @[Rob.scala 211:83 Rob.scala 211:83]
  wire  _GEN_170 = 3'h2 == dispatch_idxs_4 ? rob_info_2_busy : _GEN_169; // @[Rob.scala 211:83 Rob.scala 211:83]
  wire  _GEN_171 = 3'h3 == dispatch_idxs_4 ? rob_info_3_busy : _GEN_170; // @[Rob.scala 211:83 Rob.scala 211:83]
  wire  _GEN_172 = 3'h4 == dispatch_idxs_4 ? rob_info_4_busy : _GEN_171; // @[Rob.scala 211:83 Rob.scala 211:83]
  wire  _GEN_173 = 3'h5 == dispatch_idxs_4 ? rob_info_5_busy : _GEN_172; // @[Rob.scala 211:83 Rob.scala 211:83]
  wire  _GEN_174 = 3'h6 == dispatch_idxs_4 ? rob_info_6_busy : _GEN_173; // @[Rob.scala 211:83 Rob.scala 211:83]
  wire  _GEN_175 = 3'h7 == dispatch_idxs_4 ? rob_info_7_busy : _GEN_174; // @[Rob.scala 211:83 Rob.scala 211:83]
  wire  _ready_mask_T_25 = ~_GEN_175; // @[Rob.scala 211:83]
  wire  _GEN_177 = 3'h1 == dispatch_idxs_4 ? rob_info_1_is_valid : rob_info_0_is_valid; // @[Rob.scala 211:101 Rob.scala 211:101]
  wire  _GEN_178 = 3'h2 == dispatch_idxs_4 ? rob_info_2_is_valid : _GEN_177; // @[Rob.scala 211:101 Rob.scala 211:101]
  wire  _GEN_179 = 3'h3 == dispatch_idxs_4 ? rob_info_3_is_valid : _GEN_178; // @[Rob.scala 211:101 Rob.scala 211:101]
  wire  _GEN_180 = 3'h4 == dispatch_idxs_4 ? rob_info_4_is_valid : _GEN_179; // @[Rob.scala 211:101 Rob.scala 211:101]
  wire  _GEN_181 = 3'h5 == dispatch_idxs_4 ? rob_info_5_is_valid : _GEN_180; // @[Rob.scala 211:101 Rob.scala 211:101]
  wire  _GEN_182 = 3'h6 == dispatch_idxs_4 ? rob_info_6_is_valid : _GEN_181; // @[Rob.scala 211:101 Rob.scala 211:101]
  wire  _GEN_183 = 3'h7 == dispatch_idxs_4 ? rob_info_7_is_valid : _GEN_182; // @[Rob.scala 211:101 Rob.scala 211:101]
  wire  _GEN_185 = 3'h1 == dispatch_idxs_4 ? rob_info_1_op1_ready : rob_info_0_op1_ready; // @[Rob.scala 211:125 Rob.scala 211:125]
  wire  _GEN_186 = 3'h2 == dispatch_idxs_4 ? rob_info_2_op1_ready : _GEN_185; // @[Rob.scala 211:125 Rob.scala 211:125]
  wire  _GEN_187 = 3'h3 == dispatch_idxs_4 ? rob_info_3_op1_ready : _GEN_186; // @[Rob.scala 211:125 Rob.scala 211:125]
  wire  _GEN_188 = 3'h4 == dispatch_idxs_4 ? rob_info_4_op1_ready : _GEN_187; // @[Rob.scala 211:125 Rob.scala 211:125]
  wire  _GEN_189 = 3'h5 == dispatch_idxs_4 ? rob_info_5_op1_ready : _GEN_188; // @[Rob.scala 211:125 Rob.scala 211:125]
  wire  _GEN_190 = 3'h6 == dispatch_idxs_4 ? rob_info_6_op1_ready : _GEN_189; // @[Rob.scala 211:125 Rob.scala 211:125]
  wire  _GEN_191 = 3'h7 == dispatch_idxs_4 ? rob_info_7_op1_ready : _GEN_190; // @[Rob.scala 211:125 Rob.scala 211:125]
  wire  _GEN_193 = 3'h1 == dispatch_idxs_4 ? rob_info_1_op2_ready : rob_info_0_op2_ready; // @[Rob.scala 211:150 Rob.scala 211:150]
  wire  _GEN_194 = 3'h2 == dispatch_idxs_4 ? rob_info_2_op2_ready : _GEN_193; // @[Rob.scala 211:150 Rob.scala 211:150]
  wire  _GEN_195 = 3'h3 == dispatch_idxs_4 ? rob_info_3_op2_ready : _GEN_194; // @[Rob.scala 211:150 Rob.scala 211:150]
  wire  _GEN_196 = 3'h4 == dispatch_idxs_4 ? rob_info_4_op2_ready : _GEN_195; // @[Rob.scala 211:150 Rob.scala 211:150]
  wire  _GEN_197 = 3'h5 == dispatch_idxs_4 ? rob_info_5_op2_ready : _GEN_196; // @[Rob.scala 211:150 Rob.scala 211:150]
  wire  _GEN_198 = 3'h6 == dispatch_idxs_4 ? rob_info_6_op2_ready : _GEN_197; // @[Rob.scala 211:150 Rob.scala 211:150]
  wire  _GEN_199 = 3'h7 == dispatch_idxs_4 ? rob_info_7_op2_ready : _GEN_198; // @[Rob.scala 211:150 Rob.scala 211:150]
  wire  ready_mask_4 = ~_GEN_167 & ~_GEN_175 & _GEN_183 & _GEN_191 & _GEN_199; // @[Rob.scala 211:150]
  wire  _GEN_201 = 3'h1 == dispatch_idxs_5 ? rob_info_1_commit_ready : rob_info_0_commit_ready; // @[Rob.scala 211:54 Rob.scala 211:54]
  wire  _GEN_202 = 3'h2 == dispatch_idxs_5 ? rob_info_2_commit_ready : _GEN_201; // @[Rob.scala 211:54 Rob.scala 211:54]
  wire  _GEN_203 = 3'h3 == dispatch_idxs_5 ? rob_info_3_commit_ready : _GEN_202; // @[Rob.scala 211:54 Rob.scala 211:54]
  wire  _GEN_204 = 3'h4 == dispatch_idxs_5 ? rob_info_4_commit_ready : _GEN_203; // @[Rob.scala 211:54 Rob.scala 211:54]
  wire  _GEN_205 = 3'h5 == dispatch_idxs_5 ? rob_info_5_commit_ready : _GEN_204; // @[Rob.scala 211:54 Rob.scala 211:54]
  wire  _GEN_206 = 3'h6 == dispatch_idxs_5 ? rob_info_6_commit_ready : _GEN_205; // @[Rob.scala 211:54 Rob.scala 211:54]
  wire  _GEN_207 = 3'h7 == dispatch_idxs_5 ? rob_info_7_commit_ready : _GEN_206; // @[Rob.scala 211:54 Rob.scala 211:54]
  wire  _ready_mask_T_30 = ~_GEN_207; // @[Rob.scala 211:54]
  wire  _GEN_209 = 3'h1 == dispatch_idxs_5 ? rob_info_1_busy : rob_info_0_busy; // @[Rob.scala 211:83 Rob.scala 211:83]
  wire  _GEN_210 = 3'h2 == dispatch_idxs_5 ? rob_info_2_busy : _GEN_209; // @[Rob.scala 211:83 Rob.scala 211:83]
  wire  _GEN_211 = 3'h3 == dispatch_idxs_5 ? rob_info_3_busy : _GEN_210; // @[Rob.scala 211:83 Rob.scala 211:83]
  wire  _GEN_212 = 3'h4 == dispatch_idxs_5 ? rob_info_4_busy : _GEN_211; // @[Rob.scala 211:83 Rob.scala 211:83]
  wire  _GEN_213 = 3'h5 == dispatch_idxs_5 ? rob_info_5_busy : _GEN_212; // @[Rob.scala 211:83 Rob.scala 211:83]
  wire  _GEN_214 = 3'h6 == dispatch_idxs_5 ? rob_info_6_busy : _GEN_213; // @[Rob.scala 211:83 Rob.scala 211:83]
  wire  _GEN_215 = 3'h7 == dispatch_idxs_5 ? rob_info_7_busy : _GEN_214; // @[Rob.scala 211:83 Rob.scala 211:83]
  wire  _ready_mask_T_31 = ~_GEN_215; // @[Rob.scala 211:83]
  wire  _GEN_217 = 3'h1 == dispatch_idxs_5 ? rob_info_1_is_valid : rob_info_0_is_valid; // @[Rob.scala 211:101 Rob.scala 211:101]
  wire  _GEN_218 = 3'h2 == dispatch_idxs_5 ? rob_info_2_is_valid : _GEN_217; // @[Rob.scala 211:101 Rob.scala 211:101]
  wire  _GEN_219 = 3'h3 == dispatch_idxs_5 ? rob_info_3_is_valid : _GEN_218; // @[Rob.scala 211:101 Rob.scala 211:101]
  wire  _GEN_220 = 3'h4 == dispatch_idxs_5 ? rob_info_4_is_valid : _GEN_219; // @[Rob.scala 211:101 Rob.scala 211:101]
  wire  _GEN_221 = 3'h5 == dispatch_idxs_5 ? rob_info_5_is_valid : _GEN_220; // @[Rob.scala 211:101 Rob.scala 211:101]
  wire  _GEN_222 = 3'h6 == dispatch_idxs_5 ? rob_info_6_is_valid : _GEN_221; // @[Rob.scala 211:101 Rob.scala 211:101]
  wire  _GEN_223 = 3'h7 == dispatch_idxs_5 ? rob_info_7_is_valid : _GEN_222; // @[Rob.scala 211:101 Rob.scala 211:101]
  wire  _GEN_225 = 3'h1 == dispatch_idxs_5 ? rob_info_1_op1_ready : rob_info_0_op1_ready; // @[Rob.scala 211:125 Rob.scala 211:125]
  wire  _GEN_226 = 3'h2 == dispatch_idxs_5 ? rob_info_2_op1_ready : _GEN_225; // @[Rob.scala 211:125 Rob.scala 211:125]
  wire  _GEN_227 = 3'h3 == dispatch_idxs_5 ? rob_info_3_op1_ready : _GEN_226; // @[Rob.scala 211:125 Rob.scala 211:125]
  wire  _GEN_228 = 3'h4 == dispatch_idxs_5 ? rob_info_4_op1_ready : _GEN_227; // @[Rob.scala 211:125 Rob.scala 211:125]
  wire  _GEN_229 = 3'h5 == dispatch_idxs_5 ? rob_info_5_op1_ready : _GEN_228; // @[Rob.scala 211:125 Rob.scala 211:125]
  wire  _GEN_230 = 3'h6 == dispatch_idxs_5 ? rob_info_6_op1_ready : _GEN_229; // @[Rob.scala 211:125 Rob.scala 211:125]
  wire  _GEN_231 = 3'h7 == dispatch_idxs_5 ? rob_info_7_op1_ready : _GEN_230; // @[Rob.scala 211:125 Rob.scala 211:125]
  wire  _GEN_233 = 3'h1 == dispatch_idxs_5 ? rob_info_1_op2_ready : rob_info_0_op2_ready; // @[Rob.scala 211:150 Rob.scala 211:150]
  wire  _GEN_234 = 3'h2 == dispatch_idxs_5 ? rob_info_2_op2_ready : _GEN_233; // @[Rob.scala 211:150 Rob.scala 211:150]
  wire  _GEN_235 = 3'h3 == dispatch_idxs_5 ? rob_info_3_op2_ready : _GEN_234; // @[Rob.scala 211:150 Rob.scala 211:150]
  wire  _GEN_236 = 3'h4 == dispatch_idxs_5 ? rob_info_4_op2_ready : _GEN_235; // @[Rob.scala 211:150 Rob.scala 211:150]
  wire  _GEN_237 = 3'h5 == dispatch_idxs_5 ? rob_info_5_op2_ready : _GEN_236; // @[Rob.scala 211:150 Rob.scala 211:150]
  wire  _GEN_238 = 3'h6 == dispatch_idxs_5 ? rob_info_6_op2_ready : _GEN_237; // @[Rob.scala 211:150 Rob.scala 211:150]
  wire  _GEN_239 = 3'h7 == dispatch_idxs_5 ? rob_info_7_op2_ready : _GEN_238; // @[Rob.scala 211:150 Rob.scala 211:150]
  wire  ready_mask_5 = ~_GEN_207 & ~_GEN_215 & _GEN_223 & _GEN_231 & _GEN_239; // @[Rob.scala 211:150]
  wire  _GEN_241 = 3'h1 == dispatch_idxs_6 ? rob_info_1_commit_ready : rob_info_0_commit_ready; // @[Rob.scala 211:54 Rob.scala 211:54]
  wire  _GEN_242 = 3'h2 == dispatch_idxs_6 ? rob_info_2_commit_ready : _GEN_241; // @[Rob.scala 211:54 Rob.scala 211:54]
  wire  _GEN_243 = 3'h3 == dispatch_idxs_6 ? rob_info_3_commit_ready : _GEN_242; // @[Rob.scala 211:54 Rob.scala 211:54]
  wire  _GEN_244 = 3'h4 == dispatch_idxs_6 ? rob_info_4_commit_ready : _GEN_243; // @[Rob.scala 211:54 Rob.scala 211:54]
  wire  _GEN_245 = 3'h5 == dispatch_idxs_6 ? rob_info_5_commit_ready : _GEN_244; // @[Rob.scala 211:54 Rob.scala 211:54]
  wire  _GEN_246 = 3'h6 == dispatch_idxs_6 ? rob_info_6_commit_ready : _GEN_245; // @[Rob.scala 211:54 Rob.scala 211:54]
  wire  _GEN_247 = 3'h7 == dispatch_idxs_6 ? rob_info_7_commit_ready : _GEN_246; // @[Rob.scala 211:54 Rob.scala 211:54]
  wire  _ready_mask_T_36 = ~_GEN_247; // @[Rob.scala 211:54]
  wire  _GEN_249 = 3'h1 == dispatch_idxs_6 ? rob_info_1_busy : rob_info_0_busy; // @[Rob.scala 211:83 Rob.scala 211:83]
  wire  _GEN_250 = 3'h2 == dispatch_idxs_6 ? rob_info_2_busy : _GEN_249; // @[Rob.scala 211:83 Rob.scala 211:83]
  wire  _GEN_251 = 3'h3 == dispatch_idxs_6 ? rob_info_3_busy : _GEN_250; // @[Rob.scala 211:83 Rob.scala 211:83]
  wire  _GEN_252 = 3'h4 == dispatch_idxs_6 ? rob_info_4_busy : _GEN_251; // @[Rob.scala 211:83 Rob.scala 211:83]
  wire  _GEN_253 = 3'h5 == dispatch_idxs_6 ? rob_info_5_busy : _GEN_252; // @[Rob.scala 211:83 Rob.scala 211:83]
  wire  _GEN_254 = 3'h6 == dispatch_idxs_6 ? rob_info_6_busy : _GEN_253; // @[Rob.scala 211:83 Rob.scala 211:83]
  wire  _GEN_255 = 3'h7 == dispatch_idxs_6 ? rob_info_7_busy : _GEN_254; // @[Rob.scala 211:83 Rob.scala 211:83]
  wire  _ready_mask_T_37 = ~_GEN_255; // @[Rob.scala 211:83]
  wire  _GEN_257 = 3'h1 == dispatch_idxs_6 ? rob_info_1_is_valid : rob_info_0_is_valid; // @[Rob.scala 211:101 Rob.scala 211:101]
  wire  _GEN_258 = 3'h2 == dispatch_idxs_6 ? rob_info_2_is_valid : _GEN_257; // @[Rob.scala 211:101 Rob.scala 211:101]
  wire  _GEN_259 = 3'h3 == dispatch_idxs_6 ? rob_info_3_is_valid : _GEN_258; // @[Rob.scala 211:101 Rob.scala 211:101]
  wire  _GEN_260 = 3'h4 == dispatch_idxs_6 ? rob_info_4_is_valid : _GEN_259; // @[Rob.scala 211:101 Rob.scala 211:101]
  wire  _GEN_261 = 3'h5 == dispatch_idxs_6 ? rob_info_5_is_valid : _GEN_260; // @[Rob.scala 211:101 Rob.scala 211:101]
  wire  _GEN_262 = 3'h6 == dispatch_idxs_6 ? rob_info_6_is_valid : _GEN_261; // @[Rob.scala 211:101 Rob.scala 211:101]
  wire  _GEN_263 = 3'h7 == dispatch_idxs_6 ? rob_info_7_is_valid : _GEN_262; // @[Rob.scala 211:101 Rob.scala 211:101]
  wire  _GEN_265 = 3'h1 == dispatch_idxs_6 ? rob_info_1_op1_ready : rob_info_0_op1_ready; // @[Rob.scala 211:125 Rob.scala 211:125]
  wire  _GEN_266 = 3'h2 == dispatch_idxs_6 ? rob_info_2_op1_ready : _GEN_265; // @[Rob.scala 211:125 Rob.scala 211:125]
  wire  _GEN_267 = 3'h3 == dispatch_idxs_6 ? rob_info_3_op1_ready : _GEN_266; // @[Rob.scala 211:125 Rob.scala 211:125]
  wire  _GEN_268 = 3'h4 == dispatch_idxs_6 ? rob_info_4_op1_ready : _GEN_267; // @[Rob.scala 211:125 Rob.scala 211:125]
  wire  _GEN_269 = 3'h5 == dispatch_idxs_6 ? rob_info_5_op1_ready : _GEN_268; // @[Rob.scala 211:125 Rob.scala 211:125]
  wire  _GEN_270 = 3'h6 == dispatch_idxs_6 ? rob_info_6_op1_ready : _GEN_269; // @[Rob.scala 211:125 Rob.scala 211:125]
  wire  _GEN_271 = 3'h7 == dispatch_idxs_6 ? rob_info_7_op1_ready : _GEN_270; // @[Rob.scala 211:125 Rob.scala 211:125]
  wire  _GEN_273 = 3'h1 == dispatch_idxs_6 ? rob_info_1_op2_ready : rob_info_0_op2_ready; // @[Rob.scala 211:150 Rob.scala 211:150]
  wire  _GEN_274 = 3'h2 == dispatch_idxs_6 ? rob_info_2_op2_ready : _GEN_273; // @[Rob.scala 211:150 Rob.scala 211:150]
  wire  _GEN_275 = 3'h3 == dispatch_idxs_6 ? rob_info_3_op2_ready : _GEN_274; // @[Rob.scala 211:150 Rob.scala 211:150]
  wire  _GEN_276 = 3'h4 == dispatch_idxs_6 ? rob_info_4_op2_ready : _GEN_275; // @[Rob.scala 211:150 Rob.scala 211:150]
  wire  _GEN_277 = 3'h5 == dispatch_idxs_6 ? rob_info_5_op2_ready : _GEN_276; // @[Rob.scala 211:150 Rob.scala 211:150]
  wire  _GEN_278 = 3'h6 == dispatch_idxs_6 ? rob_info_6_op2_ready : _GEN_277; // @[Rob.scala 211:150 Rob.scala 211:150]
  wire  _GEN_279 = 3'h7 == dispatch_idxs_6 ? rob_info_7_op2_ready : _GEN_278; // @[Rob.scala 211:150 Rob.scala 211:150]
  wire  ready_mask_6 = ~_GEN_247 & ~_GEN_255 & _GEN_263 & _GEN_271 & _GEN_279; // @[Rob.scala 211:150]
  wire  _GEN_281 = 3'h1 == dispatch_idxs_7 ? rob_info_1_commit_ready : rob_info_0_commit_ready; // @[Rob.scala 211:54 Rob.scala 211:54]
  wire  _GEN_282 = 3'h2 == dispatch_idxs_7 ? rob_info_2_commit_ready : _GEN_281; // @[Rob.scala 211:54 Rob.scala 211:54]
  wire  _GEN_283 = 3'h3 == dispatch_idxs_7 ? rob_info_3_commit_ready : _GEN_282; // @[Rob.scala 211:54 Rob.scala 211:54]
  wire  _GEN_284 = 3'h4 == dispatch_idxs_7 ? rob_info_4_commit_ready : _GEN_283; // @[Rob.scala 211:54 Rob.scala 211:54]
  wire  _GEN_285 = 3'h5 == dispatch_idxs_7 ? rob_info_5_commit_ready : _GEN_284; // @[Rob.scala 211:54 Rob.scala 211:54]
  wire  _GEN_286 = 3'h6 == dispatch_idxs_7 ? rob_info_6_commit_ready : _GEN_285; // @[Rob.scala 211:54 Rob.scala 211:54]
  wire  _GEN_287 = 3'h7 == dispatch_idxs_7 ? rob_info_7_commit_ready : _GEN_286; // @[Rob.scala 211:54 Rob.scala 211:54]
  wire  _ready_mask_T_42 = ~_GEN_287; // @[Rob.scala 211:54]
  wire  _GEN_289 = 3'h1 == dispatch_idxs_7 ? rob_info_1_busy : rob_info_0_busy; // @[Rob.scala 211:83 Rob.scala 211:83]
  wire  _GEN_290 = 3'h2 == dispatch_idxs_7 ? rob_info_2_busy : _GEN_289; // @[Rob.scala 211:83 Rob.scala 211:83]
  wire  _GEN_291 = 3'h3 == dispatch_idxs_7 ? rob_info_3_busy : _GEN_290; // @[Rob.scala 211:83 Rob.scala 211:83]
  wire  _GEN_292 = 3'h4 == dispatch_idxs_7 ? rob_info_4_busy : _GEN_291; // @[Rob.scala 211:83 Rob.scala 211:83]
  wire  _GEN_293 = 3'h5 == dispatch_idxs_7 ? rob_info_5_busy : _GEN_292; // @[Rob.scala 211:83 Rob.scala 211:83]
  wire  _GEN_294 = 3'h6 == dispatch_idxs_7 ? rob_info_6_busy : _GEN_293; // @[Rob.scala 211:83 Rob.scala 211:83]
  wire  _GEN_295 = 3'h7 == dispatch_idxs_7 ? rob_info_7_busy : _GEN_294; // @[Rob.scala 211:83 Rob.scala 211:83]
  wire  _ready_mask_T_43 = ~_GEN_295; // @[Rob.scala 211:83]
  wire  _GEN_297 = 3'h1 == dispatch_idxs_7 ? rob_info_1_is_valid : rob_info_0_is_valid; // @[Rob.scala 211:101 Rob.scala 211:101]
  wire  _GEN_298 = 3'h2 == dispatch_idxs_7 ? rob_info_2_is_valid : _GEN_297; // @[Rob.scala 211:101 Rob.scala 211:101]
  wire  _GEN_299 = 3'h3 == dispatch_idxs_7 ? rob_info_3_is_valid : _GEN_298; // @[Rob.scala 211:101 Rob.scala 211:101]
  wire  _GEN_300 = 3'h4 == dispatch_idxs_7 ? rob_info_4_is_valid : _GEN_299; // @[Rob.scala 211:101 Rob.scala 211:101]
  wire  _GEN_301 = 3'h5 == dispatch_idxs_7 ? rob_info_5_is_valid : _GEN_300; // @[Rob.scala 211:101 Rob.scala 211:101]
  wire  _GEN_302 = 3'h6 == dispatch_idxs_7 ? rob_info_6_is_valid : _GEN_301; // @[Rob.scala 211:101 Rob.scala 211:101]
  wire  _GEN_303 = 3'h7 == dispatch_idxs_7 ? rob_info_7_is_valid : _GEN_302; // @[Rob.scala 211:101 Rob.scala 211:101]
  wire  _GEN_305 = 3'h1 == dispatch_idxs_7 ? rob_info_1_op1_ready : rob_info_0_op1_ready; // @[Rob.scala 211:125 Rob.scala 211:125]
  wire  _GEN_306 = 3'h2 == dispatch_idxs_7 ? rob_info_2_op1_ready : _GEN_305; // @[Rob.scala 211:125 Rob.scala 211:125]
  wire  _GEN_307 = 3'h3 == dispatch_idxs_7 ? rob_info_3_op1_ready : _GEN_306; // @[Rob.scala 211:125 Rob.scala 211:125]
  wire  _GEN_308 = 3'h4 == dispatch_idxs_7 ? rob_info_4_op1_ready : _GEN_307; // @[Rob.scala 211:125 Rob.scala 211:125]
  wire  _GEN_309 = 3'h5 == dispatch_idxs_7 ? rob_info_5_op1_ready : _GEN_308; // @[Rob.scala 211:125 Rob.scala 211:125]
  wire  _GEN_310 = 3'h6 == dispatch_idxs_7 ? rob_info_6_op1_ready : _GEN_309; // @[Rob.scala 211:125 Rob.scala 211:125]
  wire  _GEN_311 = 3'h7 == dispatch_idxs_7 ? rob_info_7_op1_ready : _GEN_310; // @[Rob.scala 211:125 Rob.scala 211:125]
  wire  _GEN_313 = 3'h1 == dispatch_idxs_7 ? rob_info_1_op2_ready : rob_info_0_op2_ready; // @[Rob.scala 211:150 Rob.scala 211:150]
  wire  _GEN_314 = 3'h2 == dispatch_idxs_7 ? rob_info_2_op2_ready : _GEN_313; // @[Rob.scala 211:150 Rob.scala 211:150]
  wire  _GEN_315 = 3'h3 == dispatch_idxs_7 ? rob_info_3_op2_ready : _GEN_314; // @[Rob.scala 211:150 Rob.scala 211:150]
  wire  _GEN_316 = 3'h4 == dispatch_idxs_7 ? rob_info_4_op2_ready : _GEN_315; // @[Rob.scala 211:150 Rob.scala 211:150]
  wire  _GEN_317 = 3'h5 == dispatch_idxs_7 ? rob_info_5_op2_ready : _GEN_316; // @[Rob.scala 211:150 Rob.scala 211:150]
  wire  _GEN_318 = 3'h6 == dispatch_idxs_7 ? rob_info_6_op2_ready : _GEN_317; // @[Rob.scala 211:150 Rob.scala 211:150]
  wire  _GEN_319 = 3'h7 == dispatch_idxs_7 ? rob_info_7_op2_ready : _GEN_318; // @[Rob.scala 211:150 Rob.scala 211:150]
  wire  ready_mask_7 = ~_GEN_287 & ~_GEN_295 & _GEN_303 & _GEN_311 & _GEN_319; // @[Rob.scala 211:150]
  wire [2:0] _GEN_321 = 3'h1 == dispatch_idxs_0 ? rob_info_1_unit_sel : rob_info_0_unit_sel; // @[Rob.scala 212:107 Rob.scala 212:107]
  wire [2:0] _GEN_322 = 3'h2 == dispatch_idxs_0 ? rob_info_2_unit_sel : _GEN_321; // @[Rob.scala 212:107 Rob.scala 212:107]
  wire [2:0] _GEN_323 = 3'h3 == dispatch_idxs_0 ? rob_info_3_unit_sel : _GEN_322; // @[Rob.scala 212:107 Rob.scala 212:107]
  wire [2:0] _GEN_324 = 3'h4 == dispatch_idxs_0 ? rob_info_4_unit_sel : _GEN_323; // @[Rob.scala 212:107 Rob.scala 212:107]
  wire [2:0] _GEN_325 = 3'h5 == dispatch_idxs_0 ? rob_info_5_unit_sel : _GEN_324; // @[Rob.scala 212:107 Rob.scala 212:107]
  wire [2:0] _GEN_326 = 3'h6 == dispatch_idxs_0 ? rob_info_6_unit_sel : _GEN_325; // @[Rob.scala 212:107 Rob.scala 212:107]
  wire [2:0] _GEN_327 = 3'h7 == dispatch_idxs_0 ? rob_info_7_unit_sel : _GEN_326; // @[Rob.scala 212:107 Rob.scala 212:107]
  wire  alu0_mask_0 = _GEN_327 == 3'h1 & ready_mask_0; // @[Rob.scala 212:126]
  wire [2:0] _GEN_329 = 3'h1 == dispatch_idxs_1 ? rob_info_1_unit_sel : rob_info_0_unit_sel; // @[Rob.scala 212:107 Rob.scala 212:107]
  wire [2:0] _GEN_330 = 3'h2 == dispatch_idxs_1 ? rob_info_2_unit_sel : _GEN_329; // @[Rob.scala 212:107 Rob.scala 212:107]
  wire [2:0] _GEN_331 = 3'h3 == dispatch_idxs_1 ? rob_info_3_unit_sel : _GEN_330; // @[Rob.scala 212:107 Rob.scala 212:107]
  wire [2:0] _GEN_332 = 3'h4 == dispatch_idxs_1 ? rob_info_4_unit_sel : _GEN_331; // @[Rob.scala 212:107 Rob.scala 212:107]
  wire [2:0] _GEN_333 = 3'h5 == dispatch_idxs_1 ? rob_info_5_unit_sel : _GEN_332; // @[Rob.scala 212:107 Rob.scala 212:107]
  wire [2:0] _GEN_334 = 3'h6 == dispatch_idxs_1 ? rob_info_6_unit_sel : _GEN_333; // @[Rob.scala 212:107 Rob.scala 212:107]
  wire [2:0] _GEN_335 = 3'h7 == dispatch_idxs_1 ? rob_info_7_unit_sel : _GEN_334; // @[Rob.scala 212:107 Rob.scala 212:107]
  wire  alu0_mask_1 = _GEN_335 == 3'h1 & ready_mask_1; // @[Rob.scala 212:126]
  wire [2:0] _GEN_337 = 3'h1 == dispatch_idxs_2 ? rob_info_1_unit_sel : rob_info_0_unit_sel; // @[Rob.scala 212:107 Rob.scala 212:107]
  wire [2:0] _GEN_338 = 3'h2 == dispatch_idxs_2 ? rob_info_2_unit_sel : _GEN_337; // @[Rob.scala 212:107 Rob.scala 212:107]
  wire [2:0] _GEN_339 = 3'h3 == dispatch_idxs_2 ? rob_info_3_unit_sel : _GEN_338; // @[Rob.scala 212:107 Rob.scala 212:107]
  wire [2:0] _GEN_340 = 3'h4 == dispatch_idxs_2 ? rob_info_4_unit_sel : _GEN_339; // @[Rob.scala 212:107 Rob.scala 212:107]
  wire [2:0] _GEN_341 = 3'h5 == dispatch_idxs_2 ? rob_info_5_unit_sel : _GEN_340; // @[Rob.scala 212:107 Rob.scala 212:107]
  wire [2:0] _GEN_342 = 3'h6 == dispatch_idxs_2 ? rob_info_6_unit_sel : _GEN_341; // @[Rob.scala 212:107 Rob.scala 212:107]
  wire [2:0] _GEN_343 = 3'h7 == dispatch_idxs_2 ? rob_info_7_unit_sel : _GEN_342; // @[Rob.scala 212:107 Rob.scala 212:107]
  wire  alu0_mask_2 = _GEN_343 == 3'h1 & ready_mask_2; // @[Rob.scala 212:126]
  wire [2:0] _GEN_345 = 3'h1 == dispatch_idxs_3 ? rob_info_1_unit_sel : rob_info_0_unit_sel; // @[Rob.scala 212:107 Rob.scala 212:107]
  wire [2:0] _GEN_346 = 3'h2 == dispatch_idxs_3 ? rob_info_2_unit_sel : _GEN_345; // @[Rob.scala 212:107 Rob.scala 212:107]
  wire [2:0] _GEN_347 = 3'h3 == dispatch_idxs_3 ? rob_info_3_unit_sel : _GEN_346; // @[Rob.scala 212:107 Rob.scala 212:107]
  wire [2:0] _GEN_348 = 3'h4 == dispatch_idxs_3 ? rob_info_4_unit_sel : _GEN_347; // @[Rob.scala 212:107 Rob.scala 212:107]
  wire [2:0] _GEN_349 = 3'h5 == dispatch_idxs_3 ? rob_info_5_unit_sel : _GEN_348; // @[Rob.scala 212:107 Rob.scala 212:107]
  wire [2:0] _GEN_350 = 3'h6 == dispatch_idxs_3 ? rob_info_6_unit_sel : _GEN_349; // @[Rob.scala 212:107 Rob.scala 212:107]
  wire [2:0] _GEN_351 = 3'h7 == dispatch_idxs_3 ? rob_info_7_unit_sel : _GEN_350; // @[Rob.scala 212:107 Rob.scala 212:107]
  wire  alu0_mask_3 = _GEN_351 == 3'h1 & ready_mask_3; // @[Rob.scala 212:126]
  wire [2:0] _GEN_353 = 3'h1 == dispatch_idxs_4 ? rob_info_1_unit_sel : rob_info_0_unit_sel; // @[Rob.scala 212:107 Rob.scala 212:107]
  wire [2:0] _GEN_354 = 3'h2 == dispatch_idxs_4 ? rob_info_2_unit_sel : _GEN_353; // @[Rob.scala 212:107 Rob.scala 212:107]
  wire [2:0] _GEN_355 = 3'h3 == dispatch_idxs_4 ? rob_info_3_unit_sel : _GEN_354; // @[Rob.scala 212:107 Rob.scala 212:107]
  wire [2:0] _GEN_356 = 3'h4 == dispatch_idxs_4 ? rob_info_4_unit_sel : _GEN_355; // @[Rob.scala 212:107 Rob.scala 212:107]
  wire [2:0] _GEN_357 = 3'h5 == dispatch_idxs_4 ? rob_info_5_unit_sel : _GEN_356; // @[Rob.scala 212:107 Rob.scala 212:107]
  wire [2:0] _GEN_358 = 3'h6 == dispatch_idxs_4 ? rob_info_6_unit_sel : _GEN_357; // @[Rob.scala 212:107 Rob.scala 212:107]
  wire [2:0] _GEN_359 = 3'h7 == dispatch_idxs_4 ? rob_info_7_unit_sel : _GEN_358; // @[Rob.scala 212:107 Rob.scala 212:107]
  wire  alu0_mask_4 = _GEN_359 == 3'h1 & ready_mask_4; // @[Rob.scala 212:126]
  wire [2:0] _GEN_361 = 3'h1 == dispatch_idxs_5 ? rob_info_1_unit_sel : rob_info_0_unit_sel; // @[Rob.scala 212:107 Rob.scala 212:107]
  wire [2:0] _GEN_362 = 3'h2 == dispatch_idxs_5 ? rob_info_2_unit_sel : _GEN_361; // @[Rob.scala 212:107 Rob.scala 212:107]
  wire [2:0] _GEN_363 = 3'h3 == dispatch_idxs_5 ? rob_info_3_unit_sel : _GEN_362; // @[Rob.scala 212:107 Rob.scala 212:107]
  wire [2:0] _GEN_364 = 3'h4 == dispatch_idxs_5 ? rob_info_4_unit_sel : _GEN_363; // @[Rob.scala 212:107 Rob.scala 212:107]
  wire [2:0] _GEN_365 = 3'h5 == dispatch_idxs_5 ? rob_info_5_unit_sel : _GEN_364; // @[Rob.scala 212:107 Rob.scala 212:107]
  wire [2:0] _GEN_366 = 3'h6 == dispatch_idxs_5 ? rob_info_6_unit_sel : _GEN_365; // @[Rob.scala 212:107 Rob.scala 212:107]
  wire [2:0] _GEN_367 = 3'h7 == dispatch_idxs_5 ? rob_info_7_unit_sel : _GEN_366; // @[Rob.scala 212:107 Rob.scala 212:107]
  wire  alu0_mask_5 = _GEN_367 == 3'h1 & ready_mask_5; // @[Rob.scala 212:126]
  wire [2:0] _GEN_369 = 3'h1 == dispatch_idxs_6 ? rob_info_1_unit_sel : rob_info_0_unit_sel; // @[Rob.scala 212:107 Rob.scala 212:107]
  wire [2:0] _GEN_370 = 3'h2 == dispatch_idxs_6 ? rob_info_2_unit_sel : _GEN_369; // @[Rob.scala 212:107 Rob.scala 212:107]
  wire [2:0] _GEN_371 = 3'h3 == dispatch_idxs_6 ? rob_info_3_unit_sel : _GEN_370; // @[Rob.scala 212:107 Rob.scala 212:107]
  wire [2:0] _GEN_372 = 3'h4 == dispatch_idxs_6 ? rob_info_4_unit_sel : _GEN_371; // @[Rob.scala 212:107 Rob.scala 212:107]
  wire [2:0] _GEN_373 = 3'h5 == dispatch_idxs_6 ? rob_info_5_unit_sel : _GEN_372; // @[Rob.scala 212:107 Rob.scala 212:107]
  wire [2:0] _GEN_374 = 3'h6 == dispatch_idxs_6 ? rob_info_6_unit_sel : _GEN_373; // @[Rob.scala 212:107 Rob.scala 212:107]
  wire [2:0] _GEN_375 = 3'h7 == dispatch_idxs_6 ? rob_info_7_unit_sel : _GEN_374; // @[Rob.scala 212:107 Rob.scala 212:107]
  wire  alu0_mask_6 = _GEN_375 == 3'h1 & ready_mask_6; // @[Rob.scala 212:126]
  wire [2:0] _GEN_377 = 3'h1 == dispatch_idxs_7 ? rob_info_1_unit_sel : rob_info_0_unit_sel; // @[Rob.scala 212:107 Rob.scala 212:107]
  wire [2:0] _GEN_378 = 3'h2 == dispatch_idxs_7 ? rob_info_2_unit_sel : _GEN_377; // @[Rob.scala 212:107 Rob.scala 212:107]
  wire [2:0] _GEN_379 = 3'h3 == dispatch_idxs_7 ? rob_info_3_unit_sel : _GEN_378; // @[Rob.scala 212:107 Rob.scala 212:107]
  wire [2:0] _GEN_380 = 3'h4 == dispatch_idxs_7 ? rob_info_4_unit_sel : _GEN_379; // @[Rob.scala 212:107 Rob.scala 212:107]
  wire [2:0] _GEN_381 = 3'h5 == dispatch_idxs_7 ? rob_info_5_unit_sel : _GEN_380; // @[Rob.scala 212:107 Rob.scala 212:107]
  wire [2:0] _GEN_382 = 3'h6 == dispatch_idxs_7 ? rob_info_6_unit_sel : _GEN_381; // @[Rob.scala 212:107 Rob.scala 212:107]
  wire [2:0] _GEN_383 = 3'h7 == dispatch_idxs_7 ? rob_info_7_unit_sel : _GEN_382; // @[Rob.scala 212:107 Rob.scala 212:107]
  wire  alu0_mask_7 = _GEN_383 == 3'h1 & ready_mask_7; // @[Rob.scala 212:126]
  wire  bju0_mask_0 = _GEN_327 == 3'h5 & ready_mask_0; // @[Rob.scala 213:127]
  wire  bju0_mask_1 = _GEN_335 == 3'h5 & ready_mask_1; // @[Rob.scala 213:127]
  wire  bju0_mask_2 = _GEN_343 == 3'h5 & ready_mask_2; // @[Rob.scala 213:127]
  wire  bju0_mask_3 = _GEN_351 == 3'h5 & ready_mask_3; // @[Rob.scala 213:127]
  wire  bju0_mask_4 = _GEN_359 == 3'h5 & ready_mask_4; // @[Rob.scala 213:127]
  wire  bju0_mask_5 = _GEN_367 == 3'h5 & ready_mask_5; // @[Rob.scala 213:127]
  wire  bju0_mask_6 = _GEN_375 == 3'h5 & ready_mask_6; // @[Rob.scala 213:127]
  wire  bju0_mask_7 = _GEN_383 == 3'h5 & ready_mask_7; // @[Rob.scala 213:127]
  wire  dispatch_mask_3_0 = _GEN_327 == 3'h4 & ready_mask_0; // @[Rob.scala 214:126]
  wire  dispatch_mask_3_1 = _GEN_335 == 3'h4 & ready_mask_1; // @[Rob.scala 214:126]
  wire  dispatch_mask_3_2 = _GEN_343 == 3'h4 & ready_mask_2; // @[Rob.scala 214:126]
  wire  dispatch_mask_3_3 = _GEN_351 == 3'h4 & ready_mask_3; // @[Rob.scala 214:126]
  wire  dispatch_mask_3_4 = _GEN_359 == 3'h4 & ready_mask_4; // @[Rob.scala 214:126]
  wire  dispatch_mask_3_5 = _GEN_367 == 3'h4 & ready_mask_5; // @[Rob.scala 214:126]
  wire  dispatch_mask_3_6 = _GEN_375 == 3'h4 & ready_mask_6; // @[Rob.scala 214:126]
  wire  dispatch_mask_3_7 = _GEN_383 == 3'h4 & ready_mask_7; // @[Rob.scala 214:126]
  wire  dispatch_mask_4_0 = _GEN_327 == 3'h3 & _ready_mask_T & _ready_mask_T_1 & _GEN_23; // @[Rob.scala 215:172]
  wire  dispatch_mask_4_1 = _GEN_335 == 3'h3 & _ready_mask_T_6 & _ready_mask_T_7 & _GEN_63; // @[Rob.scala 215:172]
  wire  dispatch_mask_4_2 = _GEN_343 == 3'h3 & _ready_mask_T_12 & _ready_mask_T_13 & _GEN_103; // @[Rob.scala 215:172]
  wire  dispatch_mask_4_3 = _GEN_351 == 3'h3 & _ready_mask_T_18 & _ready_mask_T_19 & _GEN_143; // @[Rob.scala 215:172]
  wire  dispatch_mask_4_4 = _GEN_359 == 3'h3 & _ready_mask_T_24 & _ready_mask_T_25 & _GEN_183; // @[Rob.scala 215:172]
  wire  dispatch_mask_4_5 = _GEN_367 == 3'h3 & _ready_mask_T_30 & _ready_mask_T_31 & _GEN_223; // @[Rob.scala 215:172]
  wire  dispatch_mask_4_6 = _GEN_375 == 3'h3 & _ready_mask_T_36 & _ready_mask_T_37 & _GEN_263; // @[Rob.scala 215:172]
  wire  dispatch_mask_4_7 = _GEN_383 == 3'h3 & _ready_mask_T_42 & _ready_mask_T_43 & _GEN_303; // @[Rob.scala 215:172]
  wire [7:0] _alu1_mask_enc_T = alu0_mask_7 ? 8'h80 : 8'h0; // @[Mux.scala 47:69]
  wire [7:0] _alu1_mask_enc_T_1 = alu0_mask_6 ? 8'h40 : _alu1_mask_enc_T; // @[Mux.scala 47:69]
  wire [7:0] _alu1_mask_enc_T_2 = alu0_mask_5 ? 8'h20 : _alu1_mask_enc_T_1; // @[Mux.scala 47:69]
  wire [7:0] _alu1_mask_enc_T_3 = alu0_mask_4 ? 8'h10 : _alu1_mask_enc_T_2; // @[Mux.scala 47:69]
  wire [7:0] _alu1_mask_enc_T_4 = alu0_mask_3 ? 8'h8 : _alu1_mask_enc_T_3; // @[Mux.scala 47:69]
  wire [7:0] _alu1_mask_enc_T_5 = alu0_mask_2 ? 8'h4 : _alu1_mask_enc_T_4; // @[Mux.scala 47:69]
  wire [7:0] _alu1_mask_enc_T_6 = alu0_mask_1 ? 8'h2 : _alu1_mask_enc_T_5; // @[Mux.scala 47:69]
  wire [7:0] alu1_mask_enc = alu0_mask_0 ? 8'h1 : _alu1_mask_enc_T_6; // @[Mux.scala 47:69]
  wire  alu1_mask_0 = ~alu1_mask_enc[0] & alu0_mask_0; // @[Rob.scala 217:92]
  wire  alu1_mask_1 = ~alu1_mask_enc[1] & alu0_mask_1; // @[Rob.scala 217:92]
  wire  alu1_mask_2 = ~alu1_mask_enc[2] & alu0_mask_2; // @[Rob.scala 217:92]
  wire  alu1_mask_3 = ~alu1_mask_enc[3] & alu0_mask_3; // @[Rob.scala 217:92]
  wire  alu1_mask_4 = ~alu1_mask_enc[4] & alu0_mask_4; // @[Rob.scala 217:92]
  wire  alu1_mask_5 = ~alu1_mask_enc[5] & alu0_mask_5; // @[Rob.scala 217:92]
  wire  alu1_mask_6 = ~alu1_mask_enc[6] & alu0_mask_6; // @[Rob.scala 217:92]
  wire  alu1_mask_7 = ~alu1_mask_enc[7] & alu0_mask_7; // @[Rob.scala 217:92]
  wire [2:0] _dispatch_idx_T = alu0_mask_6 ? 3'h6 : 3'h7; // @[Mux.scala 47:69]
  wire [2:0] _dispatch_idx_T_1 = alu0_mask_5 ? 3'h5 : _dispatch_idx_T; // @[Mux.scala 47:69]
  wire [2:0] _dispatch_idx_T_2 = alu0_mask_4 ? 3'h4 : _dispatch_idx_T_1; // @[Mux.scala 47:69]
  wire [2:0] _dispatch_idx_T_3 = alu0_mask_3 ? 3'h3 : _dispatch_idx_T_2; // @[Mux.scala 47:69]
  wire [2:0] _dispatch_idx_T_4 = alu0_mask_2 ? 3'h2 : _dispatch_idx_T_3; // @[Mux.scala 47:69]
  wire [2:0] _dispatch_idx_T_5 = alu0_mask_1 ? 3'h1 : _dispatch_idx_T_4; // @[Mux.scala 47:69]
  wire [2:0] dispatch_idx = alu0_mask_0 ? 3'h0 : _dispatch_idx_T_5; // @[Mux.scala 47:69]
  wire  _GEN_385 = 3'h1 == dispatch_idx ? ready_mask_1 : ready_mask_0; // @[Rob.scala 224:50 Rob.scala 224:50]
  wire  _GEN_386 = 3'h2 == dispatch_idx ? ready_mask_2 : _GEN_385; // @[Rob.scala 224:50 Rob.scala 224:50]
  wire  _GEN_387 = 3'h3 == dispatch_idx ? ready_mask_3 : _GEN_386; // @[Rob.scala 224:50 Rob.scala 224:50]
  wire  _GEN_388 = 3'h4 == dispatch_idx ? ready_mask_4 : _GEN_387; // @[Rob.scala 224:50 Rob.scala 224:50]
  wire  _GEN_389 = 3'h5 == dispatch_idx ? ready_mask_5 : _GEN_388; // @[Rob.scala 224:50 Rob.scala 224:50]
  wire  _GEN_390 = 3'h6 == dispatch_idx ? ready_mask_6 : _GEN_389; // @[Rob.scala 224:50 Rob.scala 224:50]
  wire  _GEN_391 = 3'h7 == dispatch_idx ? ready_mask_7 : _GEN_390; // @[Rob.scala 224:50 Rob.scala 224:50]
  wire  _GEN_393 = 3'h1 == dispatch_idx ? alu0_mask_1 : alu0_mask_0; // @[Rob.scala 224:50 Rob.scala 224:50]
  wire  _GEN_394 = 3'h2 == dispatch_idx ? alu0_mask_2 : _GEN_393; // @[Rob.scala 224:50 Rob.scala 224:50]
  wire  _GEN_395 = 3'h3 == dispatch_idx ? alu0_mask_3 : _GEN_394; // @[Rob.scala 224:50 Rob.scala 224:50]
  wire  _GEN_396 = 3'h4 == dispatch_idx ? alu0_mask_4 : _GEN_395; // @[Rob.scala 224:50 Rob.scala 224:50]
  wire  _GEN_397 = 3'h5 == dispatch_idx ? alu0_mask_5 : _GEN_396; // @[Rob.scala 224:50 Rob.scala 224:50]
  wire  _GEN_398 = 3'h6 == dispatch_idx ? alu0_mask_6 : _GEN_397; // @[Rob.scala 224:50 Rob.scala 224:50]
  wire  _GEN_399 = 3'h7 == dispatch_idx ? alu0_mask_7 : _GEN_398; // @[Rob.scala 224:50 Rob.scala 224:50]
  wire  dispatch_valid = _GEN_391 & _GEN_399; // @[Rob.scala 224:50]
  wire [2:0] _GEN_401 = 3'h1 == dispatch_idx ? dispatch_idxs_1 : dispatch_idxs_0; // @[Rob.scala 226:40 Rob.scala 226:40]
  wire [2:0] _GEN_402 = 3'h2 == dispatch_idx ? dispatch_idxs_2 : _GEN_401; // @[Rob.scala 226:40 Rob.scala 226:40]
  wire [2:0] _GEN_403 = 3'h3 == dispatch_idx ? dispatch_idxs_3 : _GEN_402; // @[Rob.scala 226:40 Rob.scala 226:40]
  wire [2:0] _GEN_404 = 3'h4 == dispatch_idx ? dispatch_idxs_4 : _GEN_403; // @[Rob.scala 226:40 Rob.scala 226:40]
  wire [2:0] _GEN_405 = 3'h5 == dispatch_idx ? dispatch_idxs_5 : _GEN_404; // @[Rob.scala 226:40 Rob.scala 226:40]
  wire [2:0] _GEN_406 = 3'h6 == dispatch_idx ? dispatch_idxs_6 : _GEN_405; // @[Rob.scala 226:40 Rob.scala 226:40]
  wire [2:0] _GEN_407 = 3'h7 == dispatch_idx ? dispatch_idxs_7 : _GEN_406; // @[Rob.scala 226:40 Rob.scala 226:40]
  wire [5:0] _GEN_409 = 3'h1 == _GEN_407 ? rob_info_1_uop : rob_info_0_uop; // @[Rob.scala 227:36 Rob.scala 227:36]
  wire [5:0] _GEN_410 = 3'h2 == _GEN_407 ? rob_info_2_uop : _GEN_409; // @[Rob.scala 227:36 Rob.scala 227:36]
  wire [5:0] _GEN_411 = 3'h3 == _GEN_407 ? rob_info_3_uop : _GEN_410; // @[Rob.scala 227:36 Rob.scala 227:36]
  wire [5:0] _GEN_412 = 3'h4 == _GEN_407 ? rob_info_4_uop : _GEN_411; // @[Rob.scala 227:36 Rob.scala 227:36]
  wire [5:0] _GEN_413 = 3'h5 == _GEN_407 ? rob_info_5_uop : _GEN_412; // @[Rob.scala 227:36 Rob.scala 227:36]
  wire [5:0] _GEN_414 = 3'h6 == _GEN_407 ? rob_info_6_uop : _GEN_413; // @[Rob.scala 227:36 Rob.scala 227:36]
  wire  _GEN_417 = 3'h1 == _GEN_407 ? rob_info_1_need_imm : rob_info_0_need_imm; // @[Rob.scala 228:41 Rob.scala 228:41]
  wire  _GEN_418 = 3'h2 == _GEN_407 ? rob_info_2_need_imm : _GEN_417; // @[Rob.scala 228:41 Rob.scala 228:41]
  wire  _GEN_419 = 3'h3 == _GEN_407 ? rob_info_3_need_imm : _GEN_418; // @[Rob.scala 228:41 Rob.scala 228:41]
  wire  _GEN_420 = 3'h4 == _GEN_407 ? rob_info_4_need_imm : _GEN_419; // @[Rob.scala 228:41 Rob.scala 228:41]
  wire  _GEN_421 = 3'h5 == _GEN_407 ? rob_info_5_need_imm : _GEN_420; // @[Rob.scala 228:41 Rob.scala 228:41]
  wire  _GEN_422 = 3'h6 == _GEN_407 ? rob_info_6_need_imm : _GEN_421; // @[Rob.scala 228:41 Rob.scala 228:41]
  wire [31:0] _GEN_433 = 3'h1 == _GEN_407 ? rob_info_1_op1_data : rob_info_0_op1_data; // @[Rob.scala 230:41 Rob.scala 230:41]
  wire [31:0] _GEN_434 = 3'h2 == _GEN_407 ? rob_info_2_op1_data : _GEN_433; // @[Rob.scala 230:41 Rob.scala 230:41]
  wire [31:0] _GEN_435 = 3'h3 == _GEN_407 ? rob_info_3_op1_data : _GEN_434; // @[Rob.scala 230:41 Rob.scala 230:41]
  wire [31:0] _GEN_436 = 3'h4 == _GEN_407 ? rob_info_4_op1_data : _GEN_435; // @[Rob.scala 230:41 Rob.scala 230:41]
  wire [31:0] _GEN_437 = 3'h5 == _GEN_407 ? rob_info_5_op1_data : _GEN_436; // @[Rob.scala 230:41 Rob.scala 230:41]
  wire [31:0] _GEN_438 = 3'h6 == _GEN_407 ? rob_info_6_op1_data : _GEN_437; // @[Rob.scala 230:41 Rob.scala 230:41]
  wire [31:0] _GEN_441 = 3'h1 == _GEN_407 ? rob_info_1_op2_data : rob_info_0_op2_data; // @[Rob.scala 231:41 Rob.scala 231:41]
  wire [31:0] _GEN_442 = 3'h2 == _GEN_407 ? rob_info_2_op2_data : _GEN_441; // @[Rob.scala 231:41 Rob.scala 231:41]
  wire [31:0] _GEN_443 = 3'h3 == _GEN_407 ? rob_info_3_op2_data : _GEN_442; // @[Rob.scala 231:41 Rob.scala 231:41]
  wire [31:0] _GEN_444 = 3'h4 == _GEN_407 ? rob_info_4_op2_data : _GEN_443; // @[Rob.scala 231:41 Rob.scala 231:41]
  wire [31:0] _GEN_445 = 3'h5 == _GEN_407 ? rob_info_5_op2_data : _GEN_444; // @[Rob.scala 231:41 Rob.scala 231:41]
  wire [31:0] _GEN_446 = 3'h6 == _GEN_407 ? rob_info_6_op2_data : _GEN_445; // @[Rob.scala 231:41 Rob.scala 231:41]
  wire [31:0] _GEN_449 = 3'h1 == _GEN_407 ? rob_info_1_imm_data : rob_info_0_imm_data; // @[Rob.scala 232:41 Rob.scala 232:41]
  wire [31:0] _GEN_450 = 3'h2 == _GEN_407 ? rob_info_2_imm_data : _GEN_449; // @[Rob.scala 232:41 Rob.scala 232:41]
  wire [31:0] _GEN_451 = 3'h3 == _GEN_407 ? rob_info_3_imm_data : _GEN_450; // @[Rob.scala 232:41 Rob.scala 232:41]
  wire [31:0] _GEN_452 = 3'h4 == _GEN_407 ? rob_info_4_imm_data : _GEN_451; // @[Rob.scala 232:41 Rob.scala 232:41]
  wire [31:0] _GEN_453 = 3'h5 == _GEN_407 ? rob_info_5_imm_data : _GEN_452; // @[Rob.scala 232:41 Rob.scala 232:41]
  wire [31:0] _GEN_454 = 3'h6 == _GEN_407 ? rob_info_6_imm_data : _GEN_453; // @[Rob.scala 232:41 Rob.scala 232:41]
  wire  _T_21 = ~need_flush; // @[Rob.scala 234:58]
  wire  _GEN_464 = 3'h0 == _GEN_407 | rob_info_0_busy; // @[Rob.scala 235:30 Rob.scala 235:30 Rob.scala 175:27]
  wire  _GEN_465 = 3'h1 == _GEN_407 | rob_info_1_busy; // @[Rob.scala 235:30 Rob.scala 235:30 Rob.scala 175:27]
  wire  _GEN_466 = 3'h2 == _GEN_407 | rob_info_2_busy; // @[Rob.scala 235:30 Rob.scala 235:30 Rob.scala 175:27]
  wire  _GEN_467 = 3'h3 == _GEN_407 | rob_info_3_busy; // @[Rob.scala 235:30 Rob.scala 235:30 Rob.scala 175:27]
  wire  _GEN_468 = 3'h4 == _GEN_407 | rob_info_4_busy; // @[Rob.scala 235:30 Rob.scala 235:30 Rob.scala 175:27]
  wire  _GEN_469 = 3'h5 == _GEN_407 | rob_info_5_busy; // @[Rob.scala 235:30 Rob.scala 235:30 Rob.scala 175:27]
  wire  _GEN_470 = 3'h6 == _GEN_407 | rob_info_6_busy; // @[Rob.scala 235:30 Rob.scala 235:30 Rob.scala 175:27]
  wire  _GEN_471 = 3'h7 == _GEN_407 | rob_info_7_busy; // @[Rob.scala 235:30 Rob.scala 235:30 Rob.scala 175:27]
  wire  _GEN_472 = dispatch_valid & ~need_flush ? _GEN_464 : rob_info_0_busy; // @[Rob.scala 234:71 Rob.scala 175:27]
  wire  _GEN_473 = dispatch_valid & ~need_flush ? _GEN_465 : rob_info_1_busy; // @[Rob.scala 234:71 Rob.scala 175:27]
  wire  _GEN_474 = dispatch_valid & ~need_flush ? _GEN_466 : rob_info_2_busy; // @[Rob.scala 234:71 Rob.scala 175:27]
  wire  _GEN_475 = dispatch_valid & ~need_flush ? _GEN_467 : rob_info_3_busy; // @[Rob.scala 234:71 Rob.scala 175:27]
  wire  _GEN_476 = dispatch_valid & ~need_flush ? _GEN_468 : rob_info_4_busy; // @[Rob.scala 234:71 Rob.scala 175:27]
  wire  _GEN_477 = dispatch_valid & ~need_flush ? _GEN_469 : rob_info_5_busy; // @[Rob.scala 234:71 Rob.scala 175:27]
  wire  _GEN_478 = dispatch_valid & ~need_flush ? _GEN_470 : rob_info_6_busy; // @[Rob.scala 234:71 Rob.scala 175:27]
  wire  _GEN_479 = dispatch_valid & ~need_flush ? _GEN_471 : rob_info_7_busy; // @[Rob.scala 234:71 Rob.scala 175:27]
  wire [2:0] _dispatch_idx_T_6 = alu1_mask_6 ? 3'h6 : 3'h7; // @[Mux.scala 47:69]
  wire [2:0] _dispatch_idx_T_7 = alu1_mask_5 ? 3'h5 : _dispatch_idx_T_6; // @[Mux.scala 47:69]
  wire [2:0] _dispatch_idx_T_8 = alu1_mask_4 ? 3'h4 : _dispatch_idx_T_7; // @[Mux.scala 47:69]
  wire [2:0] _dispatch_idx_T_9 = alu1_mask_3 ? 3'h3 : _dispatch_idx_T_8; // @[Mux.scala 47:69]
  wire [2:0] _dispatch_idx_T_10 = alu1_mask_2 ? 3'h2 : _dispatch_idx_T_9; // @[Mux.scala 47:69]
  wire [2:0] _dispatch_idx_T_11 = alu1_mask_1 ? 3'h1 : _dispatch_idx_T_10; // @[Mux.scala 47:69]
  wire [2:0] dispatch_idx_1 = alu1_mask_0 ? 3'h0 : _dispatch_idx_T_11; // @[Mux.scala 47:69]
  wire  _GEN_481 = 3'h1 == dispatch_idx_1 ? ready_mask_1 : ready_mask_0; // @[Rob.scala 224:50 Rob.scala 224:50]
  wire  _GEN_482 = 3'h2 == dispatch_idx_1 ? ready_mask_2 : _GEN_481; // @[Rob.scala 224:50 Rob.scala 224:50]
  wire  _GEN_483 = 3'h3 == dispatch_idx_1 ? ready_mask_3 : _GEN_482; // @[Rob.scala 224:50 Rob.scala 224:50]
  wire  _GEN_484 = 3'h4 == dispatch_idx_1 ? ready_mask_4 : _GEN_483; // @[Rob.scala 224:50 Rob.scala 224:50]
  wire  _GEN_485 = 3'h5 == dispatch_idx_1 ? ready_mask_5 : _GEN_484; // @[Rob.scala 224:50 Rob.scala 224:50]
  wire  _GEN_486 = 3'h6 == dispatch_idx_1 ? ready_mask_6 : _GEN_485; // @[Rob.scala 224:50 Rob.scala 224:50]
  wire  _GEN_487 = 3'h7 == dispatch_idx_1 ? ready_mask_7 : _GEN_486; // @[Rob.scala 224:50 Rob.scala 224:50]
  wire  _GEN_489 = 3'h1 == dispatch_idx_1 ? alu1_mask_1 : alu1_mask_0; // @[Rob.scala 224:50 Rob.scala 224:50]
  wire  _GEN_490 = 3'h2 == dispatch_idx_1 ? alu1_mask_2 : _GEN_489; // @[Rob.scala 224:50 Rob.scala 224:50]
  wire  _GEN_491 = 3'h3 == dispatch_idx_1 ? alu1_mask_3 : _GEN_490; // @[Rob.scala 224:50 Rob.scala 224:50]
  wire  _GEN_492 = 3'h4 == dispatch_idx_1 ? alu1_mask_4 : _GEN_491; // @[Rob.scala 224:50 Rob.scala 224:50]
  wire  _GEN_493 = 3'h5 == dispatch_idx_1 ? alu1_mask_5 : _GEN_492; // @[Rob.scala 224:50 Rob.scala 224:50]
  wire  _GEN_494 = 3'h6 == dispatch_idx_1 ? alu1_mask_6 : _GEN_493; // @[Rob.scala 224:50 Rob.scala 224:50]
  wire  _GEN_495 = 3'h7 == dispatch_idx_1 ? alu1_mask_7 : _GEN_494; // @[Rob.scala 224:50 Rob.scala 224:50]
  wire  dispatch_valid_1 = _GEN_487 & _GEN_495; // @[Rob.scala 224:50]
  wire [2:0] _GEN_497 = 3'h1 == dispatch_idx_1 ? dispatch_idxs_1 : dispatch_idxs_0; // @[Rob.scala 226:40 Rob.scala 226:40]
  wire [2:0] _GEN_498 = 3'h2 == dispatch_idx_1 ? dispatch_idxs_2 : _GEN_497; // @[Rob.scala 226:40 Rob.scala 226:40]
  wire [2:0] _GEN_499 = 3'h3 == dispatch_idx_1 ? dispatch_idxs_3 : _GEN_498; // @[Rob.scala 226:40 Rob.scala 226:40]
  wire [2:0] _GEN_500 = 3'h4 == dispatch_idx_1 ? dispatch_idxs_4 : _GEN_499; // @[Rob.scala 226:40 Rob.scala 226:40]
  wire [2:0] _GEN_501 = 3'h5 == dispatch_idx_1 ? dispatch_idxs_5 : _GEN_500; // @[Rob.scala 226:40 Rob.scala 226:40]
  wire [2:0] _GEN_502 = 3'h6 == dispatch_idx_1 ? dispatch_idxs_6 : _GEN_501; // @[Rob.scala 226:40 Rob.scala 226:40]
  wire [2:0] _GEN_503 = 3'h7 == dispatch_idx_1 ? dispatch_idxs_7 : _GEN_502; // @[Rob.scala 226:40 Rob.scala 226:40]
  wire [5:0] _GEN_505 = 3'h1 == _GEN_503 ? rob_info_1_uop : rob_info_0_uop; // @[Rob.scala 227:36 Rob.scala 227:36]
  wire [5:0] _GEN_506 = 3'h2 == _GEN_503 ? rob_info_2_uop : _GEN_505; // @[Rob.scala 227:36 Rob.scala 227:36]
  wire [5:0] _GEN_507 = 3'h3 == _GEN_503 ? rob_info_3_uop : _GEN_506; // @[Rob.scala 227:36 Rob.scala 227:36]
  wire [5:0] _GEN_508 = 3'h4 == _GEN_503 ? rob_info_4_uop : _GEN_507; // @[Rob.scala 227:36 Rob.scala 227:36]
  wire [5:0] _GEN_509 = 3'h5 == _GEN_503 ? rob_info_5_uop : _GEN_508; // @[Rob.scala 227:36 Rob.scala 227:36]
  wire [5:0] _GEN_510 = 3'h6 == _GEN_503 ? rob_info_6_uop : _GEN_509; // @[Rob.scala 227:36 Rob.scala 227:36]
  wire  _GEN_513 = 3'h1 == _GEN_503 ? rob_info_1_need_imm : rob_info_0_need_imm; // @[Rob.scala 228:41 Rob.scala 228:41]
  wire  _GEN_514 = 3'h2 == _GEN_503 ? rob_info_2_need_imm : _GEN_513; // @[Rob.scala 228:41 Rob.scala 228:41]
  wire  _GEN_515 = 3'h3 == _GEN_503 ? rob_info_3_need_imm : _GEN_514; // @[Rob.scala 228:41 Rob.scala 228:41]
  wire  _GEN_516 = 3'h4 == _GEN_503 ? rob_info_4_need_imm : _GEN_515; // @[Rob.scala 228:41 Rob.scala 228:41]
  wire  _GEN_517 = 3'h5 == _GEN_503 ? rob_info_5_need_imm : _GEN_516; // @[Rob.scala 228:41 Rob.scala 228:41]
  wire  _GEN_518 = 3'h6 == _GEN_503 ? rob_info_6_need_imm : _GEN_517; // @[Rob.scala 228:41 Rob.scala 228:41]
  wire [31:0] _GEN_529 = 3'h1 == _GEN_503 ? rob_info_1_op1_data : rob_info_0_op1_data; // @[Rob.scala 230:41 Rob.scala 230:41]
  wire [31:0] _GEN_530 = 3'h2 == _GEN_503 ? rob_info_2_op1_data : _GEN_529; // @[Rob.scala 230:41 Rob.scala 230:41]
  wire [31:0] _GEN_531 = 3'h3 == _GEN_503 ? rob_info_3_op1_data : _GEN_530; // @[Rob.scala 230:41 Rob.scala 230:41]
  wire [31:0] _GEN_532 = 3'h4 == _GEN_503 ? rob_info_4_op1_data : _GEN_531; // @[Rob.scala 230:41 Rob.scala 230:41]
  wire [31:0] _GEN_533 = 3'h5 == _GEN_503 ? rob_info_5_op1_data : _GEN_532; // @[Rob.scala 230:41 Rob.scala 230:41]
  wire [31:0] _GEN_534 = 3'h6 == _GEN_503 ? rob_info_6_op1_data : _GEN_533; // @[Rob.scala 230:41 Rob.scala 230:41]
  wire [31:0] _GEN_537 = 3'h1 == _GEN_503 ? rob_info_1_op2_data : rob_info_0_op2_data; // @[Rob.scala 231:41 Rob.scala 231:41]
  wire [31:0] _GEN_538 = 3'h2 == _GEN_503 ? rob_info_2_op2_data : _GEN_537; // @[Rob.scala 231:41 Rob.scala 231:41]
  wire [31:0] _GEN_539 = 3'h3 == _GEN_503 ? rob_info_3_op2_data : _GEN_538; // @[Rob.scala 231:41 Rob.scala 231:41]
  wire [31:0] _GEN_540 = 3'h4 == _GEN_503 ? rob_info_4_op2_data : _GEN_539; // @[Rob.scala 231:41 Rob.scala 231:41]
  wire [31:0] _GEN_541 = 3'h5 == _GEN_503 ? rob_info_5_op2_data : _GEN_540; // @[Rob.scala 231:41 Rob.scala 231:41]
  wire [31:0] _GEN_542 = 3'h6 == _GEN_503 ? rob_info_6_op2_data : _GEN_541; // @[Rob.scala 231:41 Rob.scala 231:41]
  wire [31:0] _GEN_545 = 3'h1 == _GEN_503 ? rob_info_1_imm_data : rob_info_0_imm_data; // @[Rob.scala 232:41 Rob.scala 232:41]
  wire [31:0] _GEN_546 = 3'h2 == _GEN_503 ? rob_info_2_imm_data : _GEN_545; // @[Rob.scala 232:41 Rob.scala 232:41]
  wire [31:0] _GEN_547 = 3'h3 == _GEN_503 ? rob_info_3_imm_data : _GEN_546; // @[Rob.scala 232:41 Rob.scala 232:41]
  wire [31:0] _GEN_548 = 3'h4 == _GEN_503 ? rob_info_4_imm_data : _GEN_547; // @[Rob.scala 232:41 Rob.scala 232:41]
  wire [31:0] _GEN_549 = 3'h5 == _GEN_503 ? rob_info_5_imm_data : _GEN_548; // @[Rob.scala 232:41 Rob.scala 232:41]
  wire [31:0] _GEN_550 = 3'h6 == _GEN_503 ? rob_info_6_imm_data : _GEN_549; // @[Rob.scala 232:41 Rob.scala 232:41]
  wire  _GEN_560 = 3'h0 == _GEN_503 | _GEN_472; // @[Rob.scala 235:30 Rob.scala 235:30]
  wire  _GEN_561 = 3'h1 == _GEN_503 | _GEN_473; // @[Rob.scala 235:30 Rob.scala 235:30]
  wire  _GEN_562 = 3'h2 == _GEN_503 | _GEN_474; // @[Rob.scala 235:30 Rob.scala 235:30]
  wire  _GEN_563 = 3'h3 == _GEN_503 | _GEN_475; // @[Rob.scala 235:30 Rob.scala 235:30]
  wire  _GEN_564 = 3'h4 == _GEN_503 | _GEN_476; // @[Rob.scala 235:30 Rob.scala 235:30]
  wire  _GEN_565 = 3'h5 == _GEN_503 | _GEN_477; // @[Rob.scala 235:30 Rob.scala 235:30]
  wire  _GEN_566 = 3'h6 == _GEN_503 | _GEN_478; // @[Rob.scala 235:30 Rob.scala 235:30]
  wire  _GEN_567 = 3'h7 == _GEN_503 | _GEN_479; // @[Rob.scala 235:30 Rob.scala 235:30]
  wire  _GEN_568 = dispatch_valid_1 & ~need_flush ? _GEN_560 : _GEN_472; // @[Rob.scala 234:71]
  wire  _GEN_569 = dispatch_valid_1 & ~need_flush ? _GEN_561 : _GEN_473; // @[Rob.scala 234:71]
  wire  _GEN_570 = dispatch_valid_1 & ~need_flush ? _GEN_562 : _GEN_474; // @[Rob.scala 234:71]
  wire  _GEN_571 = dispatch_valid_1 & ~need_flush ? _GEN_563 : _GEN_475; // @[Rob.scala 234:71]
  wire  _GEN_572 = dispatch_valid_1 & ~need_flush ? _GEN_564 : _GEN_476; // @[Rob.scala 234:71]
  wire  _GEN_573 = dispatch_valid_1 & ~need_flush ? _GEN_565 : _GEN_477; // @[Rob.scala 234:71]
  wire  _GEN_574 = dispatch_valid_1 & ~need_flush ? _GEN_566 : _GEN_478; // @[Rob.scala 234:71]
  wire  _GEN_575 = dispatch_valid_1 & ~need_flush ? _GEN_567 : _GEN_479; // @[Rob.scala 234:71]
  wire [2:0] _dispatch_idx_T_12 = bju0_mask_6 ? 3'h6 : 3'h7; // @[Mux.scala 47:69]
  wire [2:0] _dispatch_idx_T_13 = bju0_mask_5 ? 3'h5 : _dispatch_idx_T_12; // @[Mux.scala 47:69]
  wire [2:0] _dispatch_idx_T_14 = bju0_mask_4 ? 3'h4 : _dispatch_idx_T_13; // @[Mux.scala 47:69]
  wire [2:0] _dispatch_idx_T_15 = bju0_mask_3 ? 3'h3 : _dispatch_idx_T_14; // @[Mux.scala 47:69]
  wire [2:0] _dispatch_idx_T_16 = bju0_mask_2 ? 3'h2 : _dispatch_idx_T_15; // @[Mux.scala 47:69]
  wire [2:0] _dispatch_idx_T_17 = bju0_mask_1 ? 3'h1 : _dispatch_idx_T_16; // @[Mux.scala 47:69]
  wire [2:0] dispatch_idx_2 = bju0_mask_0 ? 3'h0 : _dispatch_idx_T_17; // @[Mux.scala 47:69]
  wire  _GEN_577 = 3'h1 == dispatch_idx_2 ? ready_mask_1 : ready_mask_0; // @[Rob.scala 224:50 Rob.scala 224:50]
  wire  _GEN_578 = 3'h2 == dispatch_idx_2 ? ready_mask_2 : _GEN_577; // @[Rob.scala 224:50 Rob.scala 224:50]
  wire  _GEN_579 = 3'h3 == dispatch_idx_2 ? ready_mask_3 : _GEN_578; // @[Rob.scala 224:50 Rob.scala 224:50]
  wire  _GEN_580 = 3'h4 == dispatch_idx_2 ? ready_mask_4 : _GEN_579; // @[Rob.scala 224:50 Rob.scala 224:50]
  wire  _GEN_581 = 3'h5 == dispatch_idx_2 ? ready_mask_5 : _GEN_580; // @[Rob.scala 224:50 Rob.scala 224:50]
  wire  _GEN_582 = 3'h6 == dispatch_idx_2 ? ready_mask_6 : _GEN_581; // @[Rob.scala 224:50 Rob.scala 224:50]
  wire  _GEN_583 = 3'h7 == dispatch_idx_2 ? ready_mask_7 : _GEN_582; // @[Rob.scala 224:50 Rob.scala 224:50]
  wire  _GEN_585 = 3'h1 == dispatch_idx_2 ? bju0_mask_1 : bju0_mask_0; // @[Rob.scala 224:50 Rob.scala 224:50]
  wire  _GEN_586 = 3'h2 == dispatch_idx_2 ? bju0_mask_2 : _GEN_585; // @[Rob.scala 224:50 Rob.scala 224:50]
  wire  _GEN_587 = 3'h3 == dispatch_idx_2 ? bju0_mask_3 : _GEN_586; // @[Rob.scala 224:50 Rob.scala 224:50]
  wire  _GEN_588 = 3'h4 == dispatch_idx_2 ? bju0_mask_4 : _GEN_587; // @[Rob.scala 224:50 Rob.scala 224:50]
  wire  _GEN_589 = 3'h5 == dispatch_idx_2 ? bju0_mask_5 : _GEN_588; // @[Rob.scala 224:50 Rob.scala 224:50]
  wire  _GEN_590 = 3'h6 == dispatch_idx_2 ? bju0_mask_6 : _GEN_589; // @[Rob.scala 224:50 Rob.scala 224:50]
  wire  _GEN_591 = 3'h7 == dispatch_idx_2 ? bju0_mask_7 : _GEN_590; // @[Rob.scala 224:50 Rob.scala 224:50]
  wire  dispatch_valid_2 = _GEN_583 & _GEN_591; // @[Rob.scala 224:50]
  wire [2:0] _GEN_593 = 3'h1 == dispatch_idx_2 ? dispatch_idxs_1 : dispatch_idxs_0; // @[Rob.scala 226:40 Rob.scala 226:40]
  wire [2:0] _GEN_594 = 3'h2 == dispatch_idx_2 ? dispatch_idxs_2 : _GEN_593; // @[Rob.scala 226:40 Rob.scala 226:40]
  wire [2:0] _GEN_595 = 3'h3 == dispatch_idx_2 ? dispatch_idxs_3 : _GEN_594; // @[Rob.scala 226:40 Rob.scala 226:40]
  wire [2:0] _GEN_596 = 3'h4 == dispatch_idx_2 ? dispatch_idxs_4 : _GEN_595; // @[Rob.scala 226:40 Rob.scala 226:40]
  wire [2:0] _GEN_597 = 3'h5 == dispatch_idx_2 ? dispatch_idxs_5 : _GEN_596; // @[Rob.scala 226:40 Rob.scala 226:40]
  wire [2:0] _GEN_598 = 3'h6 == dispatch_idx_2 ? dispatch_idxs_6 : _GEN_597; // @[Rob.scala 226:40 Rob.scala 226:40]
  wire [2:0] _GEN_599 = 3'h7 == dispatch_idx_2 ? dispatch_idxs_7 : _GEN_598; // @[Rob.scala 226:40 Rob.scala 226:40]
  wire [5:0] _GEN_601 = 3'h1 == _GEN_599 ? rob_info_1_uop : rob_info_0_uop; // @[Rob.scala 227:36 Rob.scala 227:36]
  wire [5:0] _GEN_602 = 3'h2 == _GEN_599 ? rob_info_2_uop : _GEN_601; // @[Rob.scala 227:36 Rob.scala 227:36]
  wire [5:0] _GEN_603 = 3'h3 == _GEN_599 ? rob_info_3_uop : _GEN_602; // @[Rob.scala 227:36 Rob.scala 227:36]
  wire [5:0] _GEN_604 = 3'h4 == _GEN_599 ? rob_info_4_uop : _GEN_603; // @[Rob.scala 227:36 Rob.scala 227:36]
  wire [5:0] _GEN_605 = 3'h5 == _GEN_599 ? rob_info_5_uop : _GEN_604; // @[Rob.scala 227:36 Rob.scala 227:36]
  wire [5:0] _GEN_606 = 3'h6 == _GEN_599 ? rob_info_6_uop : _GEN_605; // @[Rob.scala 227:36 Rob.scala 227:36]
  wire [31:0] _GEN_617 = 3'h1 == _GEN_599 ? rob_info_1_inst_addr : rob_info_0_inst_addr; // @[Rob.scala 229:42 Rob.scala 229:42]
  wire [31:0] _GEN_618 = 3'h2 == _GEN_599 ? rob_info_2_inst_addr : _GEN_617; // @[Rob.scala 229:42 Rob.scala 229:42]
  wire [31:0] _GEN_619 = 3'h3 == _GEN_599 ? rob_info_3_inst_addr : _GEN_618; // @[Rob.scala 229:42 Rob.scala 229:42]
  wire [31:0] _GEN_620 = 3'h4 == _GEN_599 ? rob_info_4_inst_addr : _GEN_619; // @[Rob.scala 229:42 Rob.scala 229:42]
  wire [31:0] _GEN_621 = 3'h5 == _GEN_599 ? rob_info_5_inst_addr : _GEN_620; // @[Rob.scala 229:42 Rob.scala 229:42]
  wire [31:0] _GEN_622 = 3'h6 == _GEN_599 ? rob_info_6_inst_addr : _GEN_621; // @[Rob.scala 229:42 Rob.scala 229:42]
  wire [31:0] _GEN_625 = 3'h1 == _GEN_599 ? rob_info_1_op1_data : rob_info_0_op1_data; // @[Rob.scala 230:41 Rob.scala 230:41]
  wire [31:0] _GEN_626 = 3'h2 == _GEN_599 ? rob_info_2_op1_data : _GEN_625; // @[Rob.scala 230:41 Rob.scala 230:41]
  wire [31:0] _GEN_627 = 3'h3 == _GEN_599 ? rob_info_3_op1_data : _GEN_626; // @[Rob.scala 230:41 Rob.scala 230:41]
  wire [31:0] _GEN_628 = 3'h4 == _GEN_599 ? rob_info_4_op1_data : _GEN_627; // @[Rob.scala 230:41 Rob.scala 230:41]
  wire [31:0] _GEN_629 = 3'h5 == _GEN_599 ? rob_info_5_op1_data : _GEN_628; // @[Rob.scala 230:41 Rob.scala 230:41]
  wire [31:0] _GEN_630 = 3'h6 == _GEN_599 ? rob_info_6_op1_data : _GEN_629; // @[Rob.scala 230:41 Rob.scala 230:41]
  wire [31:0] _GEN_633 = 3'h1 == _GEN_599 ? rob_info_1_op2_data : rob_info_0_op2_data; // @[Rob.scala 231:41 Rob.scala 231:41]
  wire [31:0] _GEN_634 = 3'h2 == _GEN_599 ? rob_info_2_op2_data : _GEN_633; // @[Rob.scala 231:41 Rob.scala 231:41]
  wire [31:0] _GEN_635 = 3'h3 == _GEN_599 ? rob_info_3_op2_data : _GEN_634; // @[Rob.scala 231:41 Rob.scala 231:41]
  wire [31:0] _GEN_636 = 3'h4 == _GEN_599 ? rob_info_4_op2_data : _GEN_635; // @[Rob.scala 231:41 Rob.scala 231:41]
  wire [31:0] _GEN_637 = 3'h5 == _GEN_599 ? rob_info_5_op2_data : _GEN_636; // @[Rob.scala 231:41 Rob.scala 231:41]
  wire [31:0] _GEN_638 = 3'h6 == _GEN_599 ? rob_info_6_op2_data : _GEN_637; // @[Rob.scala 231:41 Rob.scala 231:41]
  wire [31:0] _GEN_641 = 3'h1 == _GEN_599 ? rob_info_1_imm_data : rob_info_0_imm_data; // @[Rob.scala 232:41 Rob.scala 232:41]
  wire [31:0] _GEN_642 = 3'h2 == _GEN_599 ? rob_info_2_imm_data : _GEN_641; // @[Rob.scala 232:41 Rob.scala 232:41]
  wire [31:0] _GEN_643 = 3'h3 == _GEN_599 ? rob_info_3_imm_data : _GEN_642; // @[Rob.scala 232:41 Rob.scala 232:41]
  wire [31:0] _GEN_644 = 3'h4 == _GEN_599 ? rob_info_4_imm_data : _GEN_643; // @[Rob.scala 232:41 Rob.scala 232:41]
  wire [31:0] _GEN_645 = 3'h5 == _GEN_599 ? rob_info_5_imm_data : _GEN_644; // @[Rob.scala 232:41 Rob.scala 232:41]
  wire [31:0] _GEN_646 = 3'h6 == _GEN_599 ? rob_info_6_imm_data : _GEN_645; // @[Rob.scala 232:41 Rob.scala 232:41]
  wire  _GEN_649 = 3'h1 == _GEN_599 ? rob_info_1_predict_taken : rob_info_0_predict_taken; // @[Rob.scala 233:46 Rob.scala 233:46]
  wire  _GEN_650 = 3'h2 == _GEN_599 ? rob_info_2_predict_taken : _GEN_649; // @[Rob.scala 233:46 Rob.scala 233:46]
  wire  _GEN_651 = 3'h3 == _GEN_599 ? rob_info_3_predict_taken : _GEN_650; // @[Rob.scala 233:46 Rob.scala 233:46]
  wire  _GEN_652 = 3'h4 == _GEN_599 ? rob_info_4_predict_taken : _GEN_651; // @[Rob.scala 233:46 Rob.scala 233:46]
  wire  _GEN_653 = 3'h5 == _GEN_599 ? rob_info_5_predict_taken : _GEN_652; // @[Rob.scala 233:46 Rob.scala 233:46]
  wire  _GEN_654 = 3'h6 == _GEN_599 ? rob_info_6_predict_taken : _GEN_653; // @[Rob.scala 233:46 Rob.scala 233:46]
  wire  _GEN_656 = 3'h0 == _GEN_599 | _GEN_568; // @[Rob.scala 235:30 Rob.scala 235:30]
  wire  _GEN_657 = 3'h1 == _GEN_599 | _GEN_569; // @[Rob.scala 235:30 Rob.scala 235:30]
  wire  _GEN_658 = 3'h2 == _GEN_599 | _GEN_570; // @[Rob.scala 235:30 Rob.scala 235:30]
  wire  _GEN_659 = 3'h3 == _GEN_599 | _GEN_571; // @[Rob.scala 235:30 Rob.scala 235:30]
  wire  _GEN_660 = 3'h4 == _GEN_599 | _GEN_572; // @[Rob.scala 235:30 Rob.scala 235:30]
  wire  _GEN_661 = 3'h5 == _GEN_599 | _GEN_573; // @[Rob.scala 235:30 Rob.scala 235:30]
  wire  _GEN_662 = 3'h6 == _GEN_599 | _GEN_574; // @[Rob.scala 235:30 Rob.scala 235:30]
  wire  _GEN_663 = 3'h7 == _GEN_599 | _GEN_575; // @[Rob.scala 235:30 Rob.scala 235:30]
  wire  _GEN_664 = dispatch_valid_2 & ~need_flush ? _GEN_656 : _GEN_568; // @[Rob.scala 234:71]
  wire  _GEN_665 = dispatch_valid_2 & ~need_flush ? _GEN_657 : _GEN_569; // @[Rob.scala 234:71]
  wire  _GEN_666 = dispatch_valid_2 & ~need_flush ? _GEN_658 : _GEN_570; // @[Rob.scala 234:71]
  wire  _GEN_667 = dispatch_valid_2 & ~need_flush ? _GEN_659 : _GEN_571; // @[Rob.scala 234:71]
  wire  _GEN_668 = dispatch_valid_2 & ~need_flush ? _GEN_660 : _GEN_572; // @[Rob.scala 234:71]
  wire  _GEN_669 = dispatch_valid_2 & ~need_flush ? _GEN_661 : _GEN_573; // @[Rob.scala 234:71]
  wire  _GEN_670 = dispatch_valid_2 & ~need_flush ? _GEN_662 : _GEN_574; // @[Rob.scala 234:71]
  wire  _GEN_671 = dispatch_valid_2 & ~need_flush ? _GEN_663 : _GEN_575; // @[Rob.scala 234:71]
  wire [2:0] _dispatch_idx_T_18 = dispatch_mask_3_6 ? 3'h6 : 3'h7; // @[Mux.scala 47:69]
  wire [2:0] _dispatch_idx_T_19 = dispatch_mask_3_5 ? 3'h5 : _dispatch_idx_T_18; // @[Mux.scala 47:69]
  wire [2:0] _dispatch_idx_T_20 = dispatch_mask_3_4 ? 3'h4 : _dispatch_idx_T_19; // @[Mux.scala 47:69]
  wire [2:0] _dispatch_idx_T_21 = dispatch_mask_3_3 ? 3'h3 : _dispatch_idx_T_20; // @[Mux.scala 47:69]
  wire [2:0] _dispatch_idx_T_22 = dispatch_mask_3_2 ? 3'h2 : _dispatch_idx_T_21; // @[Mux.scala 47:69]
  wire [2:0] _dispatch_idx_T_23 = dispatch_mask_3_1 ? 3'h1 : _dispatch_idx_T_22; // @[Mux.scala 47:69]
  wire [2:0] dispatch_idx_3 = dispatch_mask_3_0 ? 3'h0 : _dispatch_idx_T_23; // @[Mux.scala 47:69]
  wire  _GEN_673 = 3'h1 == dispatch_idx_3 ? ready_mask_1 : ready_mask_0; // @[Rob.scala 224:50 Rob.scala 224:50]
  wire  _GEN_674 = 3'h2 == dispatch_idx_3 ? ready_mask_2 : _GEN_673; // @[Rob.scala 224:50 Rob.scala 224:50]
  wire  _GEN_675 = 3'h3 == dispatch_idx_3 ? ready_mask_3 : _GEN_674; // @[Rob.scala 224:50 Rob.scala 224:50]
  wire  _GEN_676 = 3'h4 == dispatch_idx_3 ? ready_mask_4 : _GEN_675; // @[Rob.scala 224:50 Rob.scala 224:50]
  wire  _GEN_677 = 3'h5 == dispatch_idx_3 ? ready_mask_5 : _GEN_676; // @[Rob.scala 224:50 Rob.scala 224:50]
  wire  _GEN_678 = 3'h6 == dispatch_idx_3 ? ready_mask_6 : _GEN_677; // @[Rob.scala 224:50 Rob.scala 224:50]
  wire  _GEN_679 = 3'h7 == dispatch_idx_3 ? ready_mask_7 : _GEN_678; // @[Rob.scala 224:50 Rob.scala 224:50]
  wire  _GEN_681 = 3'h1 == dispatch_idx_3 ? dispatch_mask_3_1 : dispatch_mask_3_0; // @[Rob.scala 224:50 Rob.scala 224:50]
  wire  _GEN_682 = 3'h2 == dispatch_idx_3 ? dispatch_mask_3_2 : _GEN_681; // @[Rob.scala 224:50 Rob.scala 224:50]
  wire  _GEN_683 = 3'h3 == dispatch_idx_3 ? dispatch_mask_3_3 : _GEN_682; // @[Rob.scala 224:50 Rob.scala 224:50]
  wire  _GEN_684 = 3'h4 == dispatch_idx_3 ? dispatch_mask_3_4 : _GEN_683; // @[Rob.scala 224:50 Rob.scala 224:50]
  wire  _GEN_685 = 3'h5 == dispatch_idx_3 ? dispatch_mask_3_5 : _GEN_684; // @[Rob.scala 224:50 Rob.scala 224:50]
  wire  _GEN_686 = 3'h6 == dispatch_idx_3 ? dispatch_mask_3_6 : _GEN_685; // @[Rob.scala 224:50 Rob.scala 224:50]
  wire  _GEN_687 = 3'h7 == dispatch_idx_3 ? dispatch_mask_3_7 : _GEN_686; // @[Rob.scala 224:50 Rob.scala 224:50]
  wire  dispatch_valid_3 = _GEN_679 & _GEN_687; // @[Rob.scala 224:50]
  wire [2:0] _GEN_689 = 3'h1 == dispatch_idx_3 ? dispatch_idxs_1 : dispatch_idxs_0; // @[Rob.scala 226:40 Rob.scala 226:40]
  wire [2:0] _GEN_690 = 3'h2 == dispatch_idx_3 ? dispatch_idxs_2 : _GEN_689; // @[Rob.scala 226:40 Rob.scala 226:40]
  wire [2:0] _GEN_691 = 3'h3 == dispatch_idx_3 ? dispatch_idxs_3 : _GEN_690; // @[Rob.scala 226:40 Rob.scala 226:40]
  wire [2:0] _GEN_692 = 3'h4 == dispatch_idx_3 ? dispatch_idxs_4 : _GEN_691; // @[Rob.scala 226:40 Rob.scala 226:40]
  wire [2:0] _GEN_693 = 3'h5 == dispatch_idx_3 ? dispatch_idxs_5 : _GEN_692; // @[Rob.scala 226:40 Rob.scala 226:40]
  wire [2:0] _GEN_694 = 3'h6 == dispatch_idx_3 ? dispatch_idxs_6 : _GEN_693; // @[Rob.scala 226:40 Rob.scala 226:40]
  wire [2:0] _GEN_695 = 3'h7 == dispatch_idx_3 ? dispatch_idxs_7 : _GEN_694; // @[Rob.scala 226:40 Rob.scala 226:40]
  wire [31:0] _GEN_721 = 3'h1 == _GEN_695 ? rob_info_1_op1_data : rob_info_0_op1_data; // @[Rob.scala 230:41 Rob.scala 230:41]
  wire [31:0] _GEN_722 = 3'h2 == _GEN_695 ? rob_info_2_op1_data : _GEN_721; // @[Rob.scala 230:41 Rob.scala 230:41]
  wire [31:0] _GEN_723 = 3'h3 == _GEN_695 ? rob_info_3_op1_data : _GEN_722; // @[Rob.scala 230:41 Rob.scala 230:41]
  wire [31:0] _GEN_724 = 3'h4 == _GEN_695 ? rob_info_4_op1_data : _GEN_723; // @[Rob.scala 230:41 Rob.scala 230:41]
  wire [31:0] _GEN_725 = 3'h5 == _GEN_695 ? rob_info_5_op1_data : _GEN_724; // @[Rob.scala 230:41 Rob.scala 230:41]
  wire [31:0] _GEN_726 = 3'h6 == _GEN_695 ? rob_info_6_op1_data : _GEN_725; // @[Rob.scala 230:41 Rob.scala 230:41]
  wire [31:0] _GEN_729 = 3'h1 == _GEN_695 ? rob_info_1_op2_data : rob_info_0_op2_data; // @[Rob.scala 231:41 Rob.scala 231:41]
  wire [31:0] _GEN_730 = 3'h2 == _GEN_695 ? rob_info_2_op2_data : _GEN_729; // @[Rob.scala 231:41 Rob.scala 231:41]
  wire [31:0] _GEN_731 = 3'h3 == _GEN_695 ? rob_info_3_op2_data : _GEN_730; // @[Rob.scala 231:41 Rob.scala 231:41]
  wire [31:0] _GEN_732 = 3'h4 == _GEN_695 ? rob_info_4_op2_data : _GEN_731; // @[Rob.scala 231:41 Rob.scala 231:41]
  wire [31:0] _GEN_733 = 3'h5 == _GEN_695 ? rob_info_5_op2_data : _GEN_732; // @[Rob.scala 231:41 Rob.scala 231:41]
  wire [31:0] _GEN_734 = 3'h6 == _GEN_695 ? rob_info_6_op2_data : _GEN_733; // @[Rob.scala 231:41 Rob.scala 231:41]
  wire  _GEN_752 = 3'h0 == _GEN_695 | _GEN_664; // @[Rob.scala 235:30 Rob.scala 235:30]
  wire  _GEN_753 = 3'h1 == _GEN_695 | _GEN_665; // @[Rob.scala 235:30 Rob.scala 235:30]
  wire  _GEN_754 = 3'h2 == _GEN_695 | _GEN_666; // @[Rob.scala 235:30 Rob.scala 235:30]
  wire  _GEN_755 = 3'h3 == _GEN_695 | _GEN_667; // @[Rob.scala 235:30 Rob.scala 235:30]
  wire  _GEN_756 = 3'h4 == _GEN_695 | _GEN_668; // @[Rob.scala 235:30 Rob.scala 235:30]
  wire  _GEN_757 = 3'h5 == _GEN_695 | _GEN_669; // @[Rob.scala 235:30 Rob.scala 235:30]
  wire  _GEN_758 = 3'h6 == _GEN_695 | _GEN_670; // @[Rob.scala 235:30 Rob.scala 235:30]
  wire  _GEN_759 = 3'h7 == _GEN_695 | _GEN_671; // @[Rob.scala 235:30 Rob.scala 235:30]
  wire  _GEN_760 = dispatch_valid_3 & ~need_flush ? _GEN_752 : _GEN_664; // @[Rob.scala 234:71]
  wire  _GEN_761 = dispatch_valid_3 & ~need_flush ? _GEN_753 : _GEN_665; // @[Rob.scala 234:71]
  wire  _GEN_762 = dispatch_valid_3 & ~need_flush ? _GEN_754 : _GEN_666; // @[Rob.scala 234:71]
  wire  _GEN_763 = dispatch_valid_3 & ~need_flush ? _GEN_755 : _GEN_667; // @[Rob.scala 234:71]
  wire  _GEN_764 = dispatch_valid_3 & ~need_flush ? _GEN_756 : _GEN_668; // @[Rob.scala 234:71]
  wire  _GEN_765 = dispatch_valid_3 & ~need_flush ? _GEN_757 : _GEN_669; // @[Rob.scala 234:71]
  wire  _GEN_766 = dispatch_valid_3 & ~need_flush ? _GEN_758 : _GEN_670; // @[Rob.scala 234:71]
  wire  _GEN_767 = dispatch_valid_3 & ~need_flush ? _GEN_759 : _GEN_671; // @[Rob.scala 234:71]
  wire [2:0] _dispatch_idx_T_24 = dispatch_mask_4_6 ? 3'h6 : 3'h7; // @[Mux.scala 47:69]
  wire [2:0] _dispatch_idx_T_25 = dispatch_mask_4_5 ? 3'h5 : _dispatch_idx_T_24; // @[Mux.scala 47:69]
  wire [2:0] _dispatch_idx_T_26 = dispatch_mask_4_4 ? 3'h4 : _dispatch_idx_T_25; // @[Mux.scala 47:69]
  wire [2:0] _dispatch_idx_T_27 = dispatch_mask_4_3 ? 3'h3 : _dispatch_idx_T_26; // @[Mux.scala 47:69]
  wire [2:0] _dispatch_idx_T_28 = dispatch_mask_4_2 ? 3'h2 : _dispatch_idx_T_27; // @[Mux.scala 47:69]
  wire [2:0] _dispatch_idx_T_29 = dispatch_mask_4_1 ? 3'h1 : _dispatch_idx_T_28; // @[Mux.scala 47:69]
  wire [2:0] dispatch_idx_4 = dispatch_mask_4_0 ? 3'h0 : _dispatch_idx_T_29; // @[Mux.scala 47:69]
  wire  _GEN_769 = 3'h1 == dispatch_idx_4 ? ready_mask_1 : ready_mask_0; // @[Rob.scala 224:50 Rob.scala 224:50]
  wire  _GEN_770 = 3'h2 == dispatch_idx_4 ? ready_mask_2 : _GEN_769; // @[Rob.scala 224:50 Rob.scala 224:50]
  wire  _GEN_771 = 3'h3 == dispatch_idx_4 ? ready_mask_3 : _GEN_770; // @[Rob.scala 224:50 Rob.scala 224:50]
  wire  _GEN_772 = 3'h4 == dispatch_idx_4 ? ready_mask_4 : _GEN_771; // @[Rob.scala 224:50 Rob.scala 224:50]
  wire  _GEN_773 = 3'h5 == dispatch_idx_4 ? ready_mask_5 : _GEN_772; // @[Rob.scala 224:50 Rob.scala 224:50]
  wire  _GEN_774 = 3'h6 == dispatch_idx_4 ? ready_mask_6 : _GEN_773; // @[Rob.scala 224:50 Rob.scala 224:50]
  wire  _GEN_775 = 3'h7 == dispatch_idx_4 ? ready_mask_7 : _GEN_774; // @[Rob.scala 224:50 Rob.scala 224:50]
  wire  _GEN_777 = 3'h1 == dispatch_idx_4 ? dispatch_mask_4_1 : dispatch_mask_4_0; // @[Rob.scala 224:50 Rob.scala 224:50]
  wire  _GEN_778 = 3'h2 == dispatch_idx_4 ? dispatch_mask_4_2 : _GEN_777; // @[Rob.scala 224:50 Rob.scala 224:50]
  wire  _GEN_779 = 3'h3 == dispatch_idx_4 ? dispatch_mask_4_3 : _GEN_778; // @[Rob.scala 224:50 Rob.scala 224:50]
  wire  _GEN_780 = 3'h4 == dispatch_idx_4 ? dispatch_mask_4_4 : _GEN_779; // @[Rob.scala 224:50 Rob.scala 224:50]
  wire  _GEN_781 = 3'h5 == dispatch_idx_4 ? dispatch_mask_4_5 : _GEN_780; // @[Rob.scala 224:50 Rob.scala 224:50]
  wire  _GEN_782 = 3'h6 == dispatch_idx_4 ? dispatch_mask_4_6 : _GEN_781; // @[Rob.scala 224:50 Rob.scala 224:50]
  wire  _GEN_783 = 3'h7 == dispatch_idx_4 ? dispatch_mask_4_7 : _GEN_782; // @[Rob.scala 224:50 Rob.scala 224:50]
  wire  dispatch_valid_4 = _GEN_775 & _GEN_783; // @[Rob.scala 224:50]
  wire [2:0] _GEN_785 = 3'h1 == dispatch_idx_4 ? dispatch_idxs_1 : dispatch_idxs_0; // @[Rob.scala 226:40 Rob.scala 226:40]
  wire [2:0] _GEN_786 = 3'h2 == dispatch_idx_4 ? dispatch_idxs_2 : _GEN_785; // @[Rob.scala 226:40 Rob.scala 226:40]
  wire [2:0] _GEN_787 = 3'h3 == dispatch_idx_4 ? dispatch_idxs_3 : _GEN_786; // @[Rob.scala 226:40 Rob.scala 226:40]
  wire [2:0] _GEN_788 = 3'h4 == dispatch_idx_4 ? dispatch_idxs_4 : _GEN_787; // @[Rob.scala 226:40 Rob.scala 226:40]
  wire [2:0] _GEN_789 = 3'h5 == dispatch_idx_4 ? dispatch_idxs_5 : _GEN_788; // @[Rob.scala 226:40 Rob.scala 226:40]
  wire [2:0] _GEN_790 = 3'h6 == dispatch_idx_4 ? dispatch_idxs_6 : _GEN_789; // @[Rob.scala 226:40 Rob.scala 226:40]
  wire [2:0] _GEN_791 = 3'h7 == dispatch_idx_4 ? dispatch_idxs_7 : _GEN_790; // @[Rob.scala 226:40 Rob.scala 226:40]
  wire [5:0] _GEN_793 = 3'h1 == _GEN_791 ? rob_info_1_uop : rob_info_0_uop; // @[Rob.scala 227:36 Rob.scala 227:36]
  wire [5:0] _GEN_794 = 3'h2 == _GEN_791 ? rob_info_2_uop : _GEN_793; // @[Rob.scala 227:36 Rob.scala 227:36]
  wire [5:0] _GEN_795 = 3'h3 == _GEN_791 ? rob_info_3_uop : _GEN_794; // @[Rob.scala 227:36 Rob.scala 227:36]
  wire [5:0] _GEN_796 = 3'h4 == _GEN_791 ? rob_info_4_uop : _GEN_795; // @[Rob.scala 227:36 Rob.scala 227:36]
  wire [5:0] _GEN_797 = 3'h5 == _GEN_791 ? rob_info_5_uop : _GEN_796; // @[Rob.scala 227:36 Rob.scala 227:36]
  wire [5:0] _GEN_798 = 3'h6 == _GEN_791 ? rob_info_6_uop : _GEN_797; // @[Rob.scala 227:36 Rob.scala 227:36]
  wire [31:0] _GEN_817 = 3'h1 == _GEN_791 ? rob_info_1_op1_data : rob_info_0_op1_data; // @[Rob.scala 230:41 Rob.scala 230:41]
  wire [31:0] _GEN_818 = 3'h2 == _GEN_791 ? rob_info_2_op1_data : _GEN_817; // @[Rob.scala 230:41 Rob.scala 230:41]
  wire [31:0] _GEN_819 = 3'h3 == _GEN_791 ? rob_info_3_op1_data : _GEN_818; // @[Rob.scala 230:41 Rob.scala 230:41]
  wire [31:0] _GEN_820 = 3'h4 == _GEN_791 ? rob_info_4_op1_data : _GEN_819; // @[Rob.scala 230:41 Rob.scala 230:41]
  wire [31:0] _GEN_821 = 3'h5 == _GEN_791 ? rob_info_5_op1_data : _GEN_820; // @[Rob.scala 230:41 Rob.scala 230:41]
  wire [31:0] _GEN_822 = 3'h6 == _GEN_791 ? rob_info_6_op1_data : _GEN_821; // @[Rob.scala 230:41 Rob.scala 230:41]
  wire [31:0] _GEN_825 = 3'h1 == _GEN_791 ? rob_info_1_op2_data : rob_info_0_op2_data; // @[Rob.scala 231:41 Rob.scala 231:41]
  wire [31:0] _GEN_826 = 3'h2 == _GEN_791 ? rob_info_2_op2_data : _GEN_825; // @[Rob.scala 231:41 Rob.scala 231:41]
  wire [31:0] _GEN_827 = 3'h3 == _GEN_791 ? rob_info_3_op2_data : _GEN_826; // @[Rob.scala 231:41 Rob.scala 231:41]
  wire [31:0] _GEN_828 = 3'h4 == _GEN_791 ? rob_info_4_op2_data : _GEN_827; // @[Rob.scala 231:41 Rob.scala 231:41]
  wire [31:0] _GEN_829 = 3'h5 == _GEN_791 ? rob_info_5_op2_data : _GEN_828; // @[Rob.scala 231:41 Rob.scala 231:41]
  wire [31:0] _GEN_830 = 3'h6 == _GEN_791 ? rob_info_6_op2_data : _GEN_829; // @[Rob.scala 231:41 Rob.scala 231:41]
  wire [31:0] _GEN_833 = 3'h1 == _GEN_791 ? rob_info_1_imm_data : rob_info_0_imm_data; // @[Rob.scala 232:41 Rob.scala 232:41]
  wire [31:0] _GEN_834 = 3'h2 == _GEN_791 ? rob_info_2_imm_data : _GEN_833; // @[Rob.scala 232:41 Rob.scala 232:41]
  wire [31:0] _GEN_835 = 3'h3 == _GEN_791 ? rob_info_3_imm_data : _GEN_834; // @[Rob.scala 232:41 Rob.scala 232:41]
  wire [31:0] _GEN_836 = 3'h4 == _GEN_791 ? rob_info_4_imm_data : _GEN_835; // @[Rob.scala 232:41 Rob.scala 232:41]
  wire [31:0] _GEN_837 = 3'h5 == _GEN_791 ? rob_info_5_imm_data : _GEN_836; // @[Rob.scala 232:41 Rob.scala 232:41]
  wire [31:0] _GEN_838 = 3'h6 == _GEN_791 ? rob_info_6_imm_data : _GEN_837; // @[Rob.scala 232:41 Rob.scala 232:41]
  wire  _GEN_848 = 3'h0 == _GEN_791 | _GEN_760; // @[Rob.scala 235:30 Rob.scala 235:30]
  wire  _GEN_849 = 3'h1 == _GEN_791 | _GEN_761; // @[Rob.scala 235:30 Rob.scala 235:30]
  wire  _GEN_850 = 3'h2 == _GEN_791 | _GEN_762; // @[Rob.scala 235:30 Rob.scala 235:30]
  wire  _GEN_851 = 3'h3 == _GEN_791 | _GEN_763; // @[Rob.scala 235:30 Rob.scala 235:30]
  wire  _GEN_852 = 3'h4 == _GEN_791 | _GEN_764; // @[Rob.scala 235:30 Rob.scala 235:30]
  wire  _GEN_853 = 3'h5 == _GEN_791 | _GEN_765; // @[Rob.scala 235:30 Rob.scala 235:30]
  wire  _GEN_854 = 3'h6 == _GEN_791 | _GEN_766; // @[Rob.scala 235:30 Rob.scala 235:30]
  wire  _GEN_855 = 3'h7 == _GEN_791 | _GEN_767; // @[Rob.scala 235:30 Rob.scala 235:30]
  wire  _GEN_856 = dispatch_valid_4 & io_dispatch_info_o_4_ready & ~need_flush ? _GEN_848 : _GEN_760; // @[Rob.scala 234:71]
  wire  _GEN_857 = dispatch_valid_4 & io_dispatch_info_o_4_ready & ~need_flush ? _GEN_849 : _GEN_761; // @[Rob.scala 234:71]
  wire  _GEN_858 = dispatch_valid_4 & io_dispatch_info_o_4_ready & ~need_flush ? _GEN_850 : _GEN_762; // @[Rob.scala 234:71]
  wire  _GEN_859 = dispatch_valid_4 & io_dispatch_info_o_4_ready & ~need_flush ? _GEN_851 : _GEN_763; // @[Rob.scala 234:71]
  wire  _GEN_860 = dispatch_valid_4 & io_dispatch_info_o_4_ready & ~need_flush ? _GEN_852 : _GEN_764; // @[Rob.scala 234:71]
  wire  _GEN_861 = dispatch_valid_4 & io_dispatch_info_o_4_ready & ~need_flush ? _GEN_853 : _GEN_765; // @[Rob.scala 234:71]
  wire  _GEN_862 = dispatch_valid_4 & io_dispatch_info_o_4_ready & ~need_flush ? _GEN_854 : _GEN_766; // @[Rob.scala 234:71]
  wire  _GEN_863 = dispatch_valid_4 & io_dispatch_info_o_4_ready & ~need_flush ? _GEN_855 : _GEN_767; // @[Rob.scala 234:71]
  wire  _GEN_864 = 3'h0 == io_rob_allocate_allocate_info_bits_0_rob_idx ? 1'h0 : rob_info_0_commit_ready; // @[Rob.scala 243:38 Rob.scala 243:38 Rob.scala 175:27]
  wire  _GEN_865 = 3'h1 == io_rob_allocate_allocate_info_bits_0_rob_idx ? 1'h0 : rob_info_1_commit_ready; // @[Rob.scala 243:38 Rob.scala 243:38 Rob.scala 175:27]
  wire  _GEN_866 = 3'h2 == io_rob_allocate_allocate_info_bits_0_rob_idx ? 1'h0 : rob_info_2_commit_ready; // @[Rob.scala 243:38 Rob.scala 243:38 Rob.scala 175:27]
  wire  _GEN_867 = 3'h3 == io_rob_allocate_allocate_info_bits_0_rob_idx ? 1'h0 : rob_info_3_commit_ready; // @[Rob.scala 243:38 Rob.scala 243:38 Rob.scala 175:27]
  wire  _GEN_868 = 3'h4 == io_rob_allocate_allocate_info_bits_0_rob_idx ? 1'h0 : rob_info_4_commit_ready; // @[Rob.scala 243:38 Rob.scala 243:38 Rob.scala 175:27]
  wire  _GEN_869 = 3'h5 == io_rob_allocate_allocate_info_bits_0_rob_idx ? 1'h0 : rob_info_5_commit_ready; // @[Rob.scala 243:38 Rob.scala 243:38 Rob.scala 175:27]
  wire  _GEN_870 = 3'h6 == io_rob_allocate_allocate_info_bits_0_rob_idx ? 1'h0 : rob_info_6_commit_ready; // @[Rob.scala 243:38 Rob.scala 243:38 Rob.scala 175:27]
  wire  _GEN_871 = 3'h7 == io_rob_allocate_allocate_info_bits_0_rob_idx ? 1'h0 : rob_info_7_commit_ready; // @[Rob.scala 243:38 Rob.scala 243:38 Rob.scala 175:27]
  wire  _GEN_872 = 3'h0 == io_rob_allocate_allocate_info_bits_0_rob_idx ? 1'h0 : _GEN_856; // @[Rob.scala 244:30 Rob.scala 244:30]
  wire  _GEN_873 = 3'h1 == io_rob_allocate_allocate_info_bits_0_rob_idx ? 1'h0 : _GEN_857; // @[Rob.scala 244:30 Rob.scala 244:30]
  wire  _GEN_874 = 3'h2 == io_rob_allocate_allocate_info_bits_0_rob_idx ? 1'h0 : _GEN_858; // @[Rob.scala 244:30 Rob.scala 244:30]
  wire  _GEN_875 = 3'h3 == io_rob_allocate_allocate_info_bits_0_rob_idx ? 1'h0 : _GEN_859; // @[Rob.scala 244:30 Rob.scala 244:30]
  wire  _GEN_876 = 3'h4 == io_rob_allocate_allocate_info_bits_0_rob_idx ? 1'h0 : _GEN_860; // @[Rob.scala 244:30 Rob.scala 244:30]
  wire  _GEN_877 = 3'h5 == io_rob_allocate_allocate_info_bits_0_rob_idx ? 1'h0 : _GEN_861; // @[Rob.scala 244:30 Rob.scala 244:30]
  wire  _GEN_878 = 3'h6 == io_rob_allocate_allocate_info_bits_0_rob_idx ? 1'h0 : _GEN_862; // @[Rob.scala 244:30 Rob.scala 244:30]
  wire  _GEN_879 = 3'h7 == io_rob_allocate_allocate_info_bits_0_rob_idx ? 1'h0 : _GEN_863; // @[Rob.scala 244:30 Rob.scala 244:30]
  wire  _GEN_880 = 3'h0 == io_rob_allocate_allocate_info_bits_0_rob_idx | rob_info_0_is_valid; // @[Rob.scala 245:34 Rob.scala 245:34 Rob.scala 175:27]
  wire  _GEN_881 = 3'h1 == io_rob_allocate_allocate_info_bits_0_rob_idx | rob_info_1_is_valid; // @[Rob.scala 245:34 Rob.scala 245:34 Rob.scala 175:27]
  wire  _GEN_882 = 3'h2 == io_rob_allocate_allocate_info_bits_0_rob_idx | rob_info_2_is_valid; // @[Rob.scala 245:34 Rob.scala 245:34 Rob.scala 175:27]
  wire  _GEN_883 = 3'h3 == io_rob_allocate_allocate_info_bits_0_rob_idx | rob_info_3_is_valid; // @[Rob.scala 245:34 Rob.scala 245:34 Rob.scala 175:27]
  wire  _GEN_884 = 3'h4 == io_rob_allocate_allocate_info_bits_0_rob_idx | rob_info_4_is_valid; // @[Rob.scala 245:34 Rob.scala 245:34 Rob.scala 175:27]
  wire  _GEN_885 = 3'h5 == io_rob_allocate_allocate_info_bits_0_rob_idx | rob_info_5_is_valid; // @[Rob.scala 245:34 Rob.scala 245:34 Rob.scala 175:27]
  wire  _GEN_886 = 3'h6 == io_rob_allocate_allocate_info_bits_0_rob_idx | rob_info_6_is_valid; // @[Rob.scala 245:34 Rob.scala 245:34 Rob.scala 175:27]
  wire  _GEN_887 = 3'h7 == io_rob_allocate_allocate_info_bits_0_rob_idx | rob_info_7_is_valid; // @[Rob.scala 245:34 Rob.scala 245:34 Rob.scala 175:27]
  wire  _GEN_888 = 3'h0 == io_rob_allocate_allocate_info_bits_0_rob_idx ? 1'h0 : rob_info_0_op1_ready; // @[Rob.scala 246:35 Rob.scala 246:35 Rob.scala 175:27]
  wire  _GEN_889 = 3'h1 == io_rob_allocate_allocate_info_bits_0_rob_idx ? 1'h0 : rob_info_1_op1_ready; // @[Rob.scala 246:35 Rob.scala 246:35 Rob.scala 175:27]
  wire  _GEN_890 = 3'h2 == io_rob_allocate_allocate_info_bits_0_rob_idx ? 1'h0 : rob_info_2_op1_ready; // @[Rob.scala 246:35 Rob.scala 246:35 Rob.scala 175:27]
  wire  _GEN_891 = 3'h3 == io_rob_allocate_allocate_info_bits_0_rob_idx ? 1'h0 : rob_info_3_op1_ready; // @[Rob.scala 246:35 Rob.scala 246:35 Rob.scala 175:27]
  wire  _GEN_892 = 3'h4 == io_rob_allocate_allocate_info_bits_0_rob_idx ? 1'h0 : rob_info_4_op1_ready; // @[Rob.scala 246:35 Rob.scala 246:35 Rob.scala 175:27]
  wire  _GEN_893 = 3'h5 == io_rob_allocate_allocate_info_bits_0_rob_idx ? 1'h0 : rob_info_5_op1_ready; // @[Rob.scala 246:35 Rob.scala 246:35 Rob.scala 175:27]
  wire  _GEN_894 = 3'h6 == io_rob_allocate_allocate_info_bits_0_rob_idx ? 1'h0 : rob_info_6_op1_ready; // @[Rob.scala 246:35 Rob.scala 246:35 Rob.scala 175:27]
  wire  _GEN_895 = 3'h7 == io_rob_allocate_allocate_info_bits_0_rob_idx ? 1'h0 : rob_info_7_op1_ready; // @[Rob.scala 246:35 Rob.scala 246:35 Rob.scala 175:27]
  wire  _GEN_896 = 3'h0 == io_rob_allocate_allocate_info_bits_0_rob_idx ? 1'h0 : rob_info_0_op2_ready; // @[Rob.scala 247:35 Rob.scala 247:35 Rob.scala 175:27]
  wire  _GEN_897 = 3'h1 == io_rob_allocate_allocate_info_bits_0_rob_idx ? 1'h0 : rob_info_1_op2_ready; // @[Rob.scala 247:35 Rob.scala 247:35 Rob.scala 175:27]
  wire  _GEN_898 = 3'h2 == io_rob_allocate_allocate_info_bits_0_rob_idx ? 1'h0 : rob_info_2_op2_ready; // @[Rob.scala 247:35 Rob.scala 247:35 Rob.scala 175:27]
  wire  _GEN_899 = 3'h3 == io_rob_allocate_allocate_info_bits_0_rob_idx ? 1'h0 : rob_info_3_op2_ready; // @[Rob.scala 247:35 Rob.scala 247:35 Rob.scala 175:27]
  wire  _GEN_900 = 3'h4 == io_rob_allocate_allocate_info_bits_0_rob_idx ? 1'h0 : rob_info_4_op2_ready; // @[Rob.scala 247:35 Rob.scala 247:35 Rob.scala 175:27]
  wire  _GEN_901 = 3'h5 == io_rob_allocate_allocate_info_bits_0_rob_idx ? 1'h0 : rob_info_5_op2_ready; // @[Rob.scala 247:35 Rob.scala 247:35 Rob.scala 175:27]
  wire  _GEN_902 = 3'h6 == io_rob_allocate_allocate_info_bits_0_rob_idx ? 1'h0 : rob_info_6_op2_ready; // @[Rob.scala 247:35 Rob.scala 247:35 Rob.scala 175:27]
  wire  _GEN_903 = 3'h7 == io_rob_allocate_allocate_info_bits_0_rob_idx ? 1'h0 : rob_info_7_op2_ready; // @[Rob.scala 247:35 Rob.scala 247:35 Rob.scala 175:27]
  wire  _GEN_904 = 3'h0 == io_rob_allocate_allocate_info_bits_0_rob_idx ? 1'h0 : rob_info_0_predict_miss; // @[Rob.scala 248:38 Rob.scala 248:38 Rob.scala 175:27]
  wire  _GEN_905 = 3'h1 == io_rob_allocate_allocate_info_bits_0_rob_idx ? 1'h0 : rob_info_1_predict_miss; // @[Rob.scala 248:38 Rob.scala 248:38 Rob.scala 175:27]
  wire  _GEN_906 = 3'h2 == io_rob_allocate_allocate_info_bits_0_rob_idx ? 1'h0 : rob_info_2_predict_miss; // @[Rob.scala 248:38 Rob.scala 248:38 Rob.scala 175:27]
  wire  _GEN_907 = 3'h3 == io_rob_allocate_allocate_info_bits_0_rob_idx ? 1'h0 : rob_info_3_predict_miss; // @[Rob.scala 248:38 Rob.scala 248:38 Rob.scala 175:27]
  wire  _GEN_908 = 3'h4 == io_rob_allocate_allocate_info_bits_0_rob_idx ? 1'h0 : rob_info_4_predict_miss; // @[Rob.scala 248:38 Rob.scala 248:38 Rob.scala 175:27]
  wire  _GEN_909 = 3'h5 == io_rob_allocate_allocate_info_bits_0_rob_idx ? 1'h0 : rob_info_5_predict_miss; // @[Rob.scala 248:38 Rob.scala 248:38 Rob.scala 175:27]
  wire  _GEN_910 = 3'h6 == io_rob_allocate_allocate_info_bits_0_rob_idx ? 1'h0 : rob_info_6_predict_miss; // @[Rob.scala 248:38 Rob.scala 248:38 Rob.scala 175:27]
  wire  _GEN_911 = 3'h7 == io_rob_allocate_allocate_info_bits_0_rob_idx ? 1'h0 : rob_info_7_predict_miss; // @[Rob.scala 248:38 Rob.scala 248:38 Rob.scala 175:27]
  wire  _GEN_912 = 3'h0 == io_rob_allocate_allocate_info_bits_0_rob_idx ? 1'h0 : rob_info_0_is_taken; // @[Rob.scala 249:34 Rob.scala 249:34 Rob.scala 175:27]
  wire  _GEN_913 = 3'h1 == io_rob_allocate_allocate_info_bits_0_rob_idx ? 1'h0 : rob_info_1_is_taken; // @[Rob.scala 249:34 Rob.scala 249:34 Rob.scala 175:27]
  wire  _GEN_914 = 3'h2 == io_rob_allocate_allocate_info_bits_0_rob_idx ? 1'h0 : rob_info_2_is_taken; // @[Rob.scala 249:34 Rob.scala 249:34 Rob.scala 175:27]
  wire  _GEN_915 = 3'h3 == io_rob_allocate_allocate_info_bits_0_rob_idx ? 1'h0 : rob_info_3_is_taken; // @[Rob.scala 249:34 Rob.scala 249:34 Rob.scala 175:27]
  wire  _GEN_916 = 3'h4 == io_rob_allocate_allocate_info_bits_0_rob_idx ? 1'h0 : rob_info_4_is_taken; // @[Rob.scala 249:34 Rob.scala 249:34 Rob.scala 175:27]
  wire  _GEN_917 = 3'h5 == io_rob_allocate_allocate_info_bits_0_rob_idx ? 1'h0 : rob_info_5_is_taken; // @[Rob.scala 249:34 Rob.scala 249:34 Rob.scala 175:27]
  wire  _GEN_918 = 3'h6 == io_rob_allocate_allocate_info_bits_0_rob_idx ? 1'h0 : rob_info_6_is_taken; // @[Rob.scala 249:34 Rob.scala 249:34 Rob.scala 175:27]
  wire  _GEN_919 = 3'h7 == io_rob_allocate_allocate_info_bits_0_rob_idx ? 1'h0 : rob_info_7_is_taken; // @[Rob.scala 249:34 Rob.scala 249:34 Rob.scala 175:27]
  wire  _GEN_920 = 3'h0 == io_rob_allocate_allocate_info_bits_0_rob_idx ? 1'h0 : rob_info_0_is_init; // @[Rob.scala 250:33 Rob.scala 250:33 Rob.scala 175:27]
  wire  _GEN_921 = 3'h1 == io_rob_allocate_allocate_info_bits_0_rob_idx ? 1'h0 : rob_info_1_is_init; // @[Rob.scala 250:33 Rob.scala 250:33 Rob.scala 175:27]
  wire  _GEN_922 = 3'h2 == io_rob_allocate_allocate_info_bits_0_rob_idx ? 1'h0 : rob_info_2_is_init; // @[Rob.scala 250:33 Rob.scala 250:33 Rob.scala 175:27]
  wire  _GEN_923 = 3'h3 == io_rob_allocate_allocate_info_bits_0_rob_idx ? 1'h0 : rob_info_3_is_init; // @[Rob.scala 250:33 Rob.scala 250:33 Rob.scala 175:27]
  wire  _GEN_924 = 3'h4 == io_rob_allocate_allocate_info_bits_0_rob_idx ? 1'h0 : rob_info_4_is_init; // @[Rob.scala 250:33 Rob.scala 250:33 Rob.scala 175:27]
  wire  _GEN_925 = 3'h5 == io_rob_allocate_allocate_info_bits_0_rob_idx ? 1'h0 : rob_info_5_is_init; // @[Rob.scala 250:33 Rob.scala 250:33 Rob.scala 175:27]
  wire  _GEN_926 = 3'h6 == io_rob_allocate_allocate_info_bits_0_rob_idx ? 1'h0 : rob_info_6_is_init; // @[Rob.scala 250:33 Rob.scala 250:33 Rob.scala 175:27]
  wire  _GEN_927 = 3'h7 == io_rob_allocate_allocate_info_bits_0_rob_idx ? 1'h0 : rob_info_7_is_init; // @[Rob.scala 250:33 Rob.scala 250:33 Rob.scala 175:27]
  wire [31:0] _GEN_928 = 3'h0 == io_rob_allocate_allocate_info_bits_0_rob_idx ?
    io_rob_allocate_allocate_info_bits_0_inst_addr : rob_info_0_inst_addr; // @[Rob.scala 251:35 Rob.scala 251:35 Rob.scala 175:27]
  wire [31:0] _GEN_929 = 3'h1 == io_rob_allocate_allocate_info_bits_0_rob_idx ?
    io_rob_allocate_allocate_info_bits_0_inst_addr : rob_info_1_inst_addr; // @[Rob.scala 251:35 Rob.scala 251:35 Rob.scala 175:27]
  wire [31:0] _GEN_930 = 3'h2 == io_rob_allocate_allocate_info_bits_0_rob_idx ?
    io_rob_allocate_allocate_info_bits_0_inst_addr : rob_info_2_inst_addr; // @[Rob.scala 251:35 Rob.scala 251:35 Rob.scala 175:27]
  wire [31:0] _GEN_931 = 3'h3 == io_rob_allocate_allocate_info_bits_0_rob_idx ?
    io_rob_allocate_allocate_info_bits_0_inst_addr : rob_info_3_inst_addr; // @[Rob.scala 251:35 Rob.scala 251:35 Rob.scala 175:27]
  wire [31:0] _GEN_932 = 3'h4 == io_rob_allocate_allocate_info_bits_0_rob_idx ?
    io_rob_allocate_allocate_info_bits_0_inst_addr : rob_info_4_inst_addr; // @[Rob.scala 251:35 Rob.scala 251:35 Rob.scala 175:27]
  wire [31:0] _GEN_933 = 3'h5 == io_rob_allocate_allocate_info_bits_0_rob_idx ?
    io_rob_allocate_allocate_info_bits_0_inst_addr : rob_info_5_inst_addr; // @[Rob.scala 251:35 Rob.scala 251:35 Rob.scala 175:27]
  wire [31:0] _GEN_934 = 3'h6 == io_rob_allocate_allocate_info_bits_0_rob_idx ?
    io_rob_allocate_allocate_info_bits_0_inst_addr : rob_info_6_inst_addr; // @[Rob.scala 251:35 Rob.scala 251:35 Rob.scala 175:27]
  wire [31:0] _GEN_935 = 3'h7 == io_rob_allocate_allocate_info_bits_0_rob_idx ?
    io_rob_allocate_allocate_info_bits_0_inst_addr : rob_info_7_inst_addr; // @[Rob.scala 251:35 Rob.scala 251:35 Rob.scala 175:27]
  wire [4:0] _GEN_936 = 3'h0 == io_rob_allocate_allocate_info_bits_0_rob_idx ?
    io_rob_allocate_allocate_info_bits_0_commit_addr[4:0] : rob_info_0_commit_addr; // @[Rob.scala 252:37 Rob.scala 252:37 Rob.scala 175:27]
  wire [4:0] _GEN_937 = 3'h1 == io_rob_allocate_allocate_info_bits_0_rob_idx ?
    io_rob_allocate_allocate_info_bits_0_commit_addr[4:0] : rob_info_1_commit_addr; // @[Rob.scala 252:37 Rob.scala 252:37 Rob.scala 175:27]
  wire [4:0] _GEN_938 = 3'h2 == io_rob_allocate_allocate_info_bits_0_rob_idx ?
    io_rob_allocate_allocate_info_bits_0_commit_addr[4:0] : rob_info_2_commit_addr; // @[Rob.scala 252:37 Rob.scala 252:37 Rob.scala 175:27]
  wire [4:0] _GEN_939 = 3'h3 == io_rob_allocate_allocate_info_bits_0_rob_idx ?
    io_rob_allocate_allocate_info_bits_0_commit_addr[4:0] : rob_info_3_commit_addr; // @[Rob.scala 252:37 Rob.scala 252:37 Rob.scala 175:27]
  wire [4:0] _GEN_940 = 3'h4 == io_rob_allocate_allocate_info_bits_0_rob_idx ?
    io_rob_allocate_allocate_info_bits_0_commit_addr[4:0] : rob_info_4_commit_addr; // @[Rob.scala 252:37 Rob.scala 252:37 Rob.scala 175:27]
  wire [4:0] _GEN_941 = 3'h5 == io_rob_allocate_allocate_info_bits_0_rob_idx ?
    io_rob_allocate_allocate_info_bits_0_commit_addr[4:0] : rob_info_5_commit_addr; // @[Rob.scala 252:37 Rob.scala 252:37 Rob.scala 175:27]
  wire [4:0] _GEN_942 = 3'h6 == io_rob_allocate_allocate_info_bits_0_rob_idx ?
    io_rob_allocate_allocate_info_bits_0_commit_addr[4:0] : rob_info_6_commit_addr; // @[Rob.scala 252:37 Rob.scala 252:37 Rob.scala 175:27]
  wire [4:0] _GEN_943 = 3'h7 == io_rob_allocate_allocate_info_bits_0_rob_idx ?
    io_rob_allocate_allocate_info_bits_0_commit_addr[4:0] : rob_info_7_commit_addr; // @[Rob.scala 252:37 Rob.scala 252:37 Rob.scala 175:27]
  wire  _GEN_960 = 3'h0 == io_rob_allocate_allocate_info_bits_0_rob_idx ? io_rob_allocate_allocate_info_bits_0_unit_sel
     == 3'h5 : rob_info_0_is_branch; // @[Rob.scala 255:35 Rob.scala 255:35 Rob.scala 175:27]
  wire  _GEN_961 = 3'h1 == io_rob_allocate_allocate_info_bits_0_rob_idx ? io_rob_allocate_allocate_info_bits_0_unit_sel
     == 3'h5 : rob_info_1_is_branch; // @[Rob.scala 255:35 Rob.scala 255:35 Rob.scala 175:27]
  wire  _GEN_962 = 3'h2 == io_rob_allocate_allocate_info_bits_0_rob_idx ? io_rob_allocate_allocate_info_bits_0_unit_sel
     == 3'h5 : rob_info_2_is_branch; // @[Rob.scala 255:35 Rob.scala 255:35 Rob.scala 175:27]
  wire  _GEN_963 = 3'h3 == io_rob_allocate_allocate_info_bits_0_rob_idx ? io_rob_allocate_allocate_info_bits_0_unit_sel
     == 3'h5 : rob_info_3_is_branch; // @[Rob.scala 255:35 Rob.scala 255:35 Rob.scala 175:27]
  wire  _GEN_964 = 3'h4 == io_rob_allocate_allocate_info_bits_0_rob_idx ? io_rob_allocate_allocate_info_bits_0_unit_sel
     == 3'h5 : rob_info_4_is_branch; // @[Rob.scala 255:35 Rob.scala 255:35 Rob.scala 175:27]
  wire  _GEN_965 = 3'h5 == io_rob_allocate_allocate_info_bits_0_rob_idx ? io_rob_allocate_allocate_info_bits_0_unit_sel
     == 3'h5 : rob_info_5_is_branch; // @[Rob.scala 255:35 Rob.scala 255:35 Rob.scala 175:27]
  wire  _GEN_966 = 3'h6 == io_rob_allocate_allocate_info_bits_0_rob_idx ? io_rob_allocate_allocate_info_bits_0_unit_sel
     == 3'h5 : rob_info_6_is_branch; // @[Rob.scala 255:35 Rob.scala 255:35 Rob.scala 175:27]
  wire  _GEN_967 = 3'h7 == io_rob_allocate_allocate_info_bits_0_rob_idx ? io_rob_allocate_allocate_info_bits_0_unit_sel
     == 3'h5 : rob_info_7_is_branch; // @[Rob.scala 255:35 Rob.scala 255:35 Rob.scala 175:27]
  wire [3:0] _GEN_976 = 3'h0 == io_rob_allocate_allocate_info_bits_0_rob_idx ?
    io_rob_allocate_allocate_info_bits_0_gh_info : rob_info_0_gh_info; // @[Rob.scala 257:33 Rob.scala 257:33 Rob.scala 175:27]
  wire [3:0] _GEN_977 = 3'h1 == io_rob_allocate_allocate_info_bits_0_rob_idx ?
    io_rob_allocate_allocate_info_bits_0_gh_info : rob_info_1_gh_info; // @[Rob.scala 257:33 Rob.scala 257:33 Rob.scala 175:27]
  wire [3:0] _GEN_978 = 3'h2 == io_rob_allocate_allocate_info_bits_0_rob_idx ?
    io_rob_allocate_allocate_info_bits_0_gh_info : rob_info_2_gh_info; // @[Rob.scala 257:33 Rob.scala 257:33 Rob.scala 175:27]
  wire [3:0] _GEN_979 = 3'h3 == io_rob_allocate_allocate_info_bits_0_rob_idx ?
    io_rob_allocate_allocate_info_bits_0_gh_info : rob_info_3_gh_info; // @[Rob.scala 257:33 Rob.scala 257:33 Rob.scala 175:27]
  wire [3:0] _GEN_980 = 3'h4 == io_rob_allocate_allocate_info_bits_0_rob_idx ?
    io_rob_allocate_allocate_info_bits_0_gh_info : rob_info_4_gh_info; // @[Rob.scala 257:33 Rob.scala 257:33 Rob.scala 175:27]
  wire [3:0] _GEN_981 = 3'h5 == io_rob_allocate_allocate_info_bits_0_rob_idx ?
    io_rob_allocate_allocate_info_bits_0_gh_info : rob_info_5_gh_info; // @[Rob.scala 257:33 Rob.scala 257:33 Rob.scala 175:27]
  wire [3:0] _GEN_982 = 3'h6 == io_rob_allocate_allocate_info_bits_0_rob_idx ?
    io_rob_allocate_allocate_info_bits_0_gh_info : rob_info_6_gh_info; // @[Rob.scala 257:33 Rob.scala 257:33 Rob.scala 175:27]
  wire [3:0] _GEN_983 = 3'h7 == io_rob_allocate_allocate_info_bits_0_rob_idx ?
    io_rob_allocate_allocate_info_bits_0_gh_info : rob_info_7_gh_info; // @[Rob.scala 257:33 Rob.scala 257:33 Rob.scala 175:27]
  wire [5:0] _GEN_984 = 3'h0 == io_rob_allocate_allocate_info_bits_0_rob_idx ? io_rob_allocate_allocate_info_bits_0_uop
     : rob_info_0_uop; // @[Rob.scala 258:29 Rob.scala 258:29 Rob.scala 175:27]
  wire [5:0] _GEN_985 = 3'h1 == io_rob_allocate_allocate_info_bits_0_rob_idx ? io_rob_allocate_allocate_info_bits_0_uop
     : rob_info_1_uop; // @[Rob.scala 258:29 Rob.scala 258:29 Rob.scala 175:27]
  wire [5:0] _GEN_986 = 3'h2 == io_rob_allocate_allocate_info_bits_0_rob_idx ? io_rob_allocate_allocate_info_bits_0_uop
     : rob_info_2_uop; // @[Rob.scala 258:29 Rob.scala 258:29 Rob.scala 175:27]
  wire [5:0] _GEN_987 = 3'h3 == io_rob_allocate_allocate_info_bits_0_rob_idx ? io_rob_allocate_allocate_info_bits_0_uop
     : rob_info_3_uop; // @[Rob.scala 258:29 Rob.scala 258:29 Rob.scala 175:27]
  wire [5:0] _GEN_988 = 3'h4 == io_rob_allocate_allocate_info_bits_0_rob_idx ? io_rob_allocate_allocate_info_bits_0_uop
     : rob_info_4_uop; // @[Rob.scala 258:29 Rob.scala 258:29 Rob.scala 175:27]
  wire [5:0] _GEN_989 = 3'h5 == io_rob_allocate_allocate_info_bits_0_rob_idx ? io_rob_allocate_allocate_info_bits_0_uop
     : rob_info_5_uop; // @[Rob.scala 258:29 Rob.scala 258:29 Rob.scala 175:27]
  wire [5:0] _GEN_990 = 3'h6 == io_rob_allocate_allocate_info_bits_0_rob_idx ? io_rob_allocate_allocate_info_bits_0_uop
     : rob_info_6_uop; // @[Rob.scala 258:29 Rob.scala 258:29 Rob.scala 175:27]
  wire [5:0] _GEN_991 = 3'h7 == io_rob_allocate_allocate_info_bits_0_rob_idx ? io_rob_allocate_allocate_info_bits_0_uop
     : rob_info_7_uop; // @[Rob.scala 258:29 Rob.scala 258:29 Rob.scala 175:27]
  wire [2:0] _GEN_992 = 3'h0 == io_rob_allocate_allocate_info_bits_0_rob_idx ?
    io_rob_allocate_allocate_info_bits_0_unit_sel : rob_info_0_unit_sel; // @[Rob.scala 259:34 Rob.scala 259:34 Rob.scala 175:27]
  wire [2:0] _GEN_993 = 3'h1 == io_rob_allocate_allocate_info_bits_0_rob_idx ?
    io_rob_allocate_allocate_info_bits_0_unit_sel : rob_info_1_unit_sel; // @[Rob.scala 259:34 Rob.scala 259:34 Rob.scala 175:27]
  wire [2:0] _GEN_994 = 3'h2 == io_rob_allocate_allocate_info_bits_0_rob_idx ?
    io_rob_allocate_allocate_info_bits_0_unit_sel : rob_info_2_unit_sel; // @[Rob.scala 259:34 Rob.scala 259:34 Rob.scala 175:27]
  wire [2:0] _GEN_995 = 3'h3 == io_rob_allocate_allocate_info_bits_0_rob_idx ?
    io_rob_allocate_allocate_info_bits_0_unit_sel : rob_info_3_unit_sel; // @[Rob.scala 259:34 Rob.scala 259:34 Rob.scala 175:27]
  wire [2:0] _GEN_996 = 3'h4 == io_rob_allocate_allocate_info_bits_0_rob_idx ?
    io_rob_allocate_allocate_info_bits_0_unit_sel : rob_info_4_unit_sel; // @[Rob.scala 259:34 Rob.scala 259:34 Rob.scala 175:27]
  wire [2:0] _GEN_997 = 3'h5 == io_rob_allocate_allocate_info_bits_0_rob_idx ?
    io_rob_allocate_allocate_info_bits_0_unit_sel : rob_info_5_unit_sel; // @[Rob.scala 259:34 Rob.scala 259:34 Rob.scala 175:27]
  wire [2:0] _GEN_998 = 3'h6 == io_rob_allocate_allocate_info_bits_0_rob_idx ?
    io_rob_allocate_allocate_info_bits_0_unit_sel : rob_info_6_unit_sel; // @[Rob.scala 259:34 Rob.scala 259:34 Rob.scala 175:27]
  wire [2:0] _GEN_999 = 3'h7 == io_rob_allocate_allocate_info_bits_0_rob_idx ?
    io_rob_allocate_allocate_info_bits_0_unit_sel : rob_info_7_unit_sel; // @[Rob.scala 259:34 Rob.scala 259:34 Rob.scala 175:27]
  wire  _GEN_1000 = 3'h0 == io_rob_allocate_allocate_info_bits_0_rob_idx ? io_rob_allocate_allocate_info_bits_0_need_imm
     : rob_info_0_need_imm; // @[Rob.scala 260:34 Rob.scala 260:34 Rob.scala 175:27]
  wire  _GEN_1001 = 3'h1 == io_rob_allocate_allocate_info_bits_0_rob_idx ? io_rob_allocate_allocate_info_bits_0_need_imm
     : rob_info_1_need_imm; // @[Rob.scala 260:34 Rob.scala 260:34 Rob.scala 175:27]
  wire  _GEN_1002 = 3'h2 == io_rob_allocate_allocate_info_bits_0_rob_idx ? io_rob_allocate_allocate_info_bits_0_need_imm
     : rob_info_2_need_imm; // @[Rob.scala 260:34 Rob.scala 260:34 Rob.scala 175:27]
  wire  _GEN_1003 = 3'h3 == io_rob_allocate_allocate_info_bits_0_rob_idx ? io_rob_allocate_allocate_info_bits_0_need_imm
     : rob_info_3_need_imm; // @[Rob.scala 260:34 Rob.scala 260:34 Rob.scala 175:27]
  wire  _GEN_1004 = 3'h4 == io_rob_allocate_allocate_info_bits_0_rob_idx ? io_rob_allocate_allocate_info_bits_0_need_imm
     : rob_info_4_need_imm; // @[Rob.scala 260:34 Rob.scala 260:34 Rob.scala 175:27]
  wire  _GEN_1005 = 3'h5 == io_rob_allocate_allocate_info_bits_0_rob_idx ? io_rob_allocate_allocate_info_bits_0_need_imm
     : rob_info_5_need_imm; // @[Rob.scala 260:34 Rob.scala 260:34 Rob.scala 175:27]
  wire  _GEN_1006 = 3'h6 == io_rob_allocate_allocate_info_bits_0_rob_idx ? io_rob_allocate_allocate_info_bits_0_need_imm
     : rob_info_6_need_imm; // @[Rob.scala 260:34 Rob.scala 260:34 Rob.scala 175:27]
  wire  _GEN_1007 = 3'h7 == io_rob_allocate_allocate_info_bits_0_rob_idx ? io_rob_allocate_allocate_info_bits_0_need_imm
     : rob_info_7_need_imm; // @[Rob.scala 260:34 Rob.scala 260:34 Rob.scala 175:27]
  wire [31:0] _GEN_1008 = 3'h0 == io_rob_allocate_allocate_info_bits_0_rob_idx ?
    io_rob_allocate_allocate_info_bits_0_imm_data : rob_info_0_imm_data; // @[Rob.scala 261:34 Rob.scala 261:34 Rob.scala 175:27]
  wire [31:0] _GEN_1009 = 3'h1 == io_rob_allocate_allocate_info_bits_0_rob_idx ?
    io_rob_allocate_allocate_info_bits_0_imm_data : rob_info_1_imm_data; // @[Rob.scala 261:34 Rob.scala 261:34 Rob.scala 175:27]
  wire [31:0] _GEN_1010 = 3'h2 == io_rob_allocate_allocate_info_bits_0_rob_idx ?
    io_rob_allocate_allocate_info_bits_0_imm_data : rob_info_2_imm_data; // @[Rob.scala 261:34 Rob.scala 261:34 Rob.scala 175:27]
  wire [31:0] _GEN_1011 = 3'h3 == io_rob_allocate_allocate_info_bits_0_rob_idx ?
    io_rob_allocate_allocate_info_bits_0_imm_data : rob_info_3_imm_data; // @[Rob.scala 261:34 Rob.scala 261:34 Rob.scala 175:27]
  wire [31:0] _GEN_1012 = 3'h4 == io_rob_allocate_allocate_info_bits_0_rob_idx ?
    io_rob_allocate_allocate_info_bits_0_imm_data : rob_info_4_imm_data; // @[Rob.scala 261:34 Rob.scala 261:34 Rob.scala 175:27]
  wire [31:0] _GEN_1013 = 3'h5 == io_rob_allocate_allocate_info_bits_0_rob_idx ?
    io_rob_allocate_allocate_info_bits_0_imm_data : rob_info_5_imm_data; // @[Rob.scala 261:34 Rob.scala 261:34 Rob.scala 175:27]
  wire [31:0] _GEN_1014 = 3'h6 == io_rob_allocate_allocate_info_bits_0_rob_idx ?
    io_rob_allocate_allocate_info_bits_0_imm_data : rob_info_6_imm_data; // @[Rob.scala 261:34 Rob.scala 261:34 Rob.scala 175:27]
  wire [31:0] _GEN_1015 = 3'h7 == io_rob_allocate_allocate_info_bits_0_rob_idx ?
    io_rob_allocate_allocate_info_bits_0_imm_data : rob_info_7_imm_data; // @[Rob.scala 261:34 Rob.scala 261:34 Rob.scala 175:27]
  wire  _GEN_1016 = 3'h0 == io_rob_allocate_allocate_info_bits_0_rob_idx ?
    io_rob_allocate_allocate_info_bits_0_flush_on_commit : rob_info_0_flush_on_commit; // @[Rob.scala 262:41 Rob.scala 262:41 Rob.scala 175:27]
  wire  _GEN_1017 = 3'h1 == io_rob_allocate_allocate_info_bits_0_rob_idx ?
    io_rob_allocate_allocate_info_bits_0_flush_on_commit : rob_info_1_flush_on_commit; // @[Rob.scala 262:41 Rob.scala 262:41 Rob.scala 175:27]
  wire  _GEN_1018 = 3'h2 == io_rob_allocate_allocate_info_bits_0_rob_idx ?
    io_rob_allocate_allocate_info_bits_0_flush_on_commit : rob_info_2_flush_on_commit; // @[Rob.scala 262:41 Rob.scala 262:41 Rob.scala 175:27]
  wire  _GEN_1019 = 3'h3 == io_rob_allocate_allocate_info_bits_0_rob_idx ?
    io_rob_allocate_allocate_info_bits_0_flush_on_commit : rob_info_3_flush_on_commit; // @[Rob.scala 262:41 Rob.scala 262:41 Rob.scala 175:27]
  wire  _GEN_1020 = 3'h4 == io_rob_allocate_allocate_info_bits_0_rob_idx ?
    io_rob_allocate_allocate_info_bits_0_flush_on_commit : rob_info_4_flush_on_commit; // @[Rob.scala 262:41 Rob.scala 262:41 Rob.scala 175:27]
  wire  _GEN_1021 = 3'h5 == io_rob_allocate_allocate_info_bits_0_rob_idx ?
    io_rob_allocate_allocate_info_bits_0_flush_on_commit : rob_info_5_flush_on_commit; // @[Rob.scala 262:41 Rob.scala 262:41 Rob.scala 175:27]
  wire  _GEN_1022 = 3'h6 == io_rob_allocate_allocate_info_bits_0_rob_idx ?
    io_rob_allocate_allocate_info_bits_0_flush_on_commit : rob_info_6_flush_on_commit; // @[Rob.scala 262:41 Rob.scala 262:41 Rob.scala 175:27]
  wire  _GEN_1023 = 3'h7 == io_rob_allocate_allocate_info_bits_0_rob_idx ?
    io_rob_allocate_allocate_info_bits_0_flush_on_commit : rob_info_7_flush_on_commit; // @[Rob.scala 262:41 Rob.scala 262:41 Rob.scala 175:27]
  wire  _GEN_1024 = 3'h0 == io_rob_allocate_allocate_info_bits_0_rob_idx ?
    io_rob_allocate_allocate_info_bits_0_predict_taken : rob_info_0_predict_taken; // @[Rob.scala 263:39 Rob.scala 263:39 Rob.scala 175:27]
  wire  _GEN_1025 = 3'h1 == io_rob_allocate_allocate_info_bits_0_rob_idx ?
    io_rob_allocate_allocate_info_bits_0_predict_taken : rob_info_1_predict_taken; // @[Rob.scala 263:39 Rob.scala 263:39 Rob.scala 175:27]
  wire  _GEN_1026 = 3'h2 == io_rob_allocate_allocate_info_bits_0_rob_idx ?
    io_rob_allocate_allocate_info_bits_0_predict_taken : rob_info_2_predict_taken; // @[Rob.scala 263:39 Rob.scala 263:39 Rob.scala 175:27]
  wire  _GEN_1027 = 3'h3 == io_rob_allocate_allocate_info_bits_0_rob_idx ?
    io_rob_allocate_allocate_info_bits_0_predict_taken : rob_info_3_predict_taken; // @[Rob.scala 263:39 Rob.scala 263:39 Rob.scala 175:27]
  wire  _GEN_1028 = 3'h4 == io_rob_allocate_allocate_info_bits_0_rob_idx ?
    io_rob_allocate_allocate_info_bits_0_predict_taken : rob_info_4_predict_taken; // @[Rob.scala 263:39 Rob.scala 263:39 Rob.scala 175:27]
  wire  _GEN_1029 = 3'h5 == io_rob_allocate_allocate_info_bits_0_rob_idx ?
    io_rob_allocate_allocate_info_bits_0_predict_taken : rob_info_5_predict_taken; // @[Rob.scala 263:39 Rob.scala 263:39 Rob.scala 175:27]
  wire  _GEN_1030 = 3'h6 == io_rob_allocate_allocate_info_bits_0_rob_idx ?
    io_rob_allocate_allocate_info_bits_0_predict_taken : rob_info_6_predict_taken; // @[Rob.scala 263:39 Rob.scala 263:39 Rob.scala 175:27]
  wire  _GEN_1031 = 3'h7 == io_rob_allocate_allocate_info_bits_0_rob_idx ?
    io_rob_allocate_allocate_info_bits_0_predict_taken : rob_info_7_predict_taken; // @[Rob.scala 263:39 Rob.scala 263:39 Rob.scala 175:27]
  wire  _GEN_1032 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_864 : rob_info_0_commit_ready; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1033 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_865 : rob_info_1_commit_ready; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1034 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_866 : rob_info_2_commit_ready; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1035 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_867 : rob_info_3_commit_ready; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1036 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_868 : rob_info_4_commit_ready; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1037 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_869 : rob_info_5_commit_ready; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1038 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_870 : rob_info_6_commit_ready; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1039 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_871 : rob_info_7_commit_ready; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1040 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_872 : _GEN_856; // @[Rob.scala 242:112]
  wire  _GEN_1041 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_873 : _GEN_857; // @[Rob.scala 242:112]
  wire  _GEN_1042 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_874 : _GEN_858; // @[Rob.scala 242:112]
  wire  _GEN_1043 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_875 : _GEN_859; // @[Rob.scala 242:112]
  wire  _GEN_1044 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_876 : _GEN_860; // @[Rob.scala 242:112]
  wire  _GEN_1045 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_877 : _GEN_861; // @[Rob.scala 242:112]
  wire  _GEN_1046 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_878 : _GEN_862; // @[Rob.scala 242:112]
  wire  _GEN_1047 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_879 : _GEN_863; // @[Rob.scala 242:112]
  wire  _GEN_1048 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_880 : rob_info_0_is_valid; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1049 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_881 : rob_info_1_is_valid; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1050 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_882 : rob_info_2_is_valid; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1051 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_883 : rob_info_3_is_valid; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1052 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_884 : rob_info_4_is_valid; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1053 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_885 : rob_info_5_is_valid; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1054 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_886 : rob_info_6_is_valid; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1055 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_887 : rob_info_7_is_valid; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1056 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_888 : rob_info_0_op1_ready; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1057 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_889 : rob_info_1_op1_ready; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1058 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_890 : rob_info_2_op1_ready; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1059 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_891 : rob_info_3_op1_ready; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1060 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_892 : rob_info_4_op1_ready; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1061 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_893 : rob_info_5_op1_ready; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1062 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_894 : rob_info_6_op1_ready; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1063 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_895 : rob_info_7_op1_ready; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1064 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_896 : rob_info_0_op2_ready; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1065 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_897 : rob_info_1_op2_ready; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1066 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_898 : rob_info_2_op2_ready; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1067 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_899 : rob_info_3_op2_ready; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1068 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_900 : rob_info_4_op2_ready; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1069 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_901 : rob_info_5_op2_ready; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1070 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_902 : rob_info_6_op2_ready; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1071 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_903 : rob_info_7_op2_ready; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1072 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_904 : rob_info_0_predict_miss; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1073 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_905 : rob_info_1_predict_miss; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1074 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_906 : rob_info_2_predict_miss; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1075 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_907 : rob_info_3_predict_miss; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1076 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_908 : rob_info_4_predict_miss; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1077 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_909 : rob_info_5_predict_miss; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1078 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_910 : rob_info_6_predict_miss; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1079 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_911 : rob_info_7_predict_miss; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1080 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_912 : rob_info_0_is_taken; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1081 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_913 : rob_info_1_is_taken; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1082 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_914 : rob_info_2_is_taken; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1083 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_915 : rob_info_3_is_taken; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1084 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_916 : rob_info_4_is_taken; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1085 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_917 : rob_info_5_is_taken; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1086 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_918 : rob_info_6_is_taken; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1087 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_919 : rob_info_7_is_taken; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1088 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_920 : rob_info_0_is_init; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1089 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_921 : rob_info_1_is_init; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1090 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_922 : rob_info_2_is_init; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1091 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_923 : rob_info_3_is_init; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1092 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_924 : rob_info_4_is_init; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1093 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_925 : rob_info_5_is_init; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1094 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_926 : rob_info_6_is_init; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1095 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_927 : rob_info_7_is_init; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire [31:0] _GEN_1096 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21
     ? _GEN_928 : rob_info_0_inst_addr; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire [31:0] _GEN_1097 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21
     ? _GEN_929 : rob_info_1_inst_addr; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire [31:0] _GEN_1098 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21
     ? _GEN_930 : rob_info_2_inst_addr; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire [31:0] _GEN_1099 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21
     ? _GEN_931 : rob_info_3_inst_addr; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire [31:0] _GEN_1100 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21
     ? _GEN_932 : rob_info_4_inst_addr; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire [31:0] _GEN_1101 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21
     ? _GEN_933 : rob_info_5_inst_addr; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire [31:0] _GEN_1102 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21
     ? _GEN_934 : rob_info_6_inst_addr; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire [31:0] _GEN_1103 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21
     ? _GEN_935 : rob_info_7_inst_addr; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire [4:0] _GEN_1104 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21
     ? _GEN_936 : rob_info_0_commit_addr; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire [4:0] _GEN_1105 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21
     ? _GEN_937 : rob_info_1_commit_addr; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire [4:0] _GEN_1106 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21
     ? _GEN_938 : rob_info_2_commit_addr; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire [4:0] _GEN_1107 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21
     ? _GEN_939 : rob_info_3_commit_addr; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire [4:0] _GEN_1108 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21
     ? _GEN_940 : rob_info_4_commit_addr; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire [4:0] _GEN_1109 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21
     ? _GEN_941 : rob_info_5_commit_addr; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire [4:0] _GEN_1110 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21
     ? _GEN_942 : rob_info_6_commit_addr; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire [4:0] _GEN_1111 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21
     ? _GEN_943 : rob_info_7_commit_addr; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1128 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_960 : rob_info_0_is_branch; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1129 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_961 : rob_info_1_is_branch; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1130 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_962 : rob_info_2_is_branch; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1131 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_963 : rob_info_3_is_branch; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1132 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_964 : rob_info_4_is_branch; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1133 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_965 : rob_info_5_is_branch; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1134 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_966 : rob_info_6_is_branch; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1135 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_967 : rob_info_7_is_branch; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire [3:0] _GEN_1144 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21
     ? _GEN_976 : rob_info_0_gh_info; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire [3:0] _GEN_1145 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21
     ? _GEN_977 : rob_info_1_gh_info; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire [3:0] _GEN_1146 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21
     ? _GEN_978 : rob_info_2_gh_info; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire [3:0] _GEN_1147 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21
     ? _GEN_979 : rob_info_3_gh_info; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire [3:0] _GEN_1148 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21
     ? _GEN_980 : rob_info_4_gh_info; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire [3:0] _GEN_1149 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21
     ? _GEN_981 : rob_info_5_gh_info; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire [3:0] _GEN_1150 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21
     ? _GEN_982 : rob_info_6_gh_info; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire [3:0] _GEN_1151 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21
     ? _GEN_983 : rob_info_7_gh_info; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire [5:0] _GEN_1152 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21
     ? _GEN_984 : rob_info_0_uop; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire [5:0] _GEN_1153 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21
     ? _GEN_985 : rob_info_1_uop; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire [5:0] _GEN_1154 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21
     ? _GEN_986 : rob_info_2_uop; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire [5:0] _GEN_1155 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21
     ? _GEN_987 : rob_info_3_uop; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire [5:0] _GEN_1156 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21
     ? _GEN_988 : rob_info_4_uop; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire [5:0] _GEN_1157 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21
     ? _GEN_989 : rob_info_5_uop; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire [5:0] _GEN_1158 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21
     ? _GEN_990 : rob_info_6_uop; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire [5:0] _GEN_1159 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21
     ? _GEN_991 : rob_info_7_uop; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire [2:0] _GEN_1160 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21
     ? _GEN_992 : rob_info_0_unit_sel; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire [2:0] _GEN_1161 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21
     ? _GEN_993 : rob_info_1_unit_sel; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire [2:0] _GEN_1162 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21
     ? _GEN_994 : rob_info_2_unit_sel; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire [2:0] _GEN_1163 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21
     ? _GEN_995 : rob_info_3_unit_sel; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire [2:0] _GEN_1164 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21
     ? _GEN_996 : rob_info_4_unit_sel; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire [2:0] _GEN_1165 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21
     ? _GEN_997 : rob_info_5_unit_sel; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire [2:0] _GEN_1166 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21
     ? _GEN_998 : rob_info_6_unit_sel; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire [2:0] _GEN_1167 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21
     ? _GEN_999 : rob_info_7_unit_sel; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1168 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_1000 : rob_info_0_need_imm; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1169 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_1001 : rob_info_1_need_imm; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1170 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_1002 : rob_info_2_need_imm; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1171 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_1003 : rob_info_3_need_imm; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1172 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_1004 : rob_info_4_need_imm; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1173 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_1005 : rob_info_5_need_imm; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1174 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_1006 : rob_info_6_need_imm; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1175 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_1007 : rob_info_7_need_imm; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire [31:0] _GEN_1176 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21
     ? _GEN_1008 : rob_info_0_imm_data; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire [31:0] _GEN_1177 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21
     ? _GEN_1009 : rob_info_1_imm_data; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire [31:0] _GEN_1178 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21
     ? _GEN_1010 : rob_info_2_imm_data; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire [31:0] _GEN_1179 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21
     ? _GEN_1011 : rob_info_3_imm_data; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire [31:0] _GEN_1180 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21
     ? _GEN_1012 : rob_info_4_imm_data; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire [31:0] _GEN_1181 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21
     ? _GEN_1013 : rob_info_5_imm_data; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire [31:0] _GEN_1182 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21
     ? _GEN_1014 : rob_info_6_imm_data; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire [31:0] _GEN_1183 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21
     ? _GEN_1015 : rob_info_7_imm_data; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1184 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_1016 : rob_info_0_flush_on_commit; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1185 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_1017 : rob_info_1_flush_on_commit; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1186 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_1018 : rob_info_2_flush_on_commit; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1187 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_1019 : rob_info_3_flush_on_commit; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1188 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_1020 : rob_info_4_flush_on_commit; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1189 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_1021 : rob_info_5_flush_on_commit; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1190 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_1022 : rob_info_6_flush_on_commit; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1191 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_1023 : rob_info_7_flush_on_commit; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1192 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_1024 : rob_info_0_predict_taken; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1193 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_1025 : rob_info_1_predict_taken; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1194 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_1026 : rob_info_2_predict_taken; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1195 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_1027 : rob_info_3_predict_taken; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1196 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_1028 : rob_info_4_predict_taken; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1197 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_1029 : rob_info_5_predict_taken; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1198 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_1030 : rob_info_6_predict_taken; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1199 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_0_inst_valid & _T_21 ?
    _GEN_1031 : rob_info_7_predict_taken; // @[Rob.scala 242:112 Rob.scala 175:27]
  wire  _GEN_1200 = 3'h0 == io_rob_allocate_allocate_info_bits_1_rob_idx ? 1'h0 : _GEN_1032; // @[Rob.scala 243:38 Rob.scala 243:38]
  wire  _GEN_1201 = 3'h1 == io_rob_allocate_allocate_info_bits_1_rob_idx ? 1'h0 : _GEN_1033; // @[Rob.scala 243:38 Rob.scala 243:38]
  wire  _GEN_1202 = 3'h2 == io_rob_allocate_allocate_info_bits_1_rob_idx ? 1'h0 : _GEN_1034; // @[Rob.scala 243:38 Rob.scala 243:38]
  wire  _GEN_1203 = 3'h3 == io_rob_allocate_allocate_info_bits_1_rob_idx ? 1'h0 : _GEN_1035; // @[Rob.scala 243:38 Rob.scala 243:38]
  wire  _GEN_1204 = 3'h4 == io_rob_allocate_allocate_info_bits_1_rob_idx ? 1'h0 : _GEN_1036; // @[Rob.scala 243:38 Rob.scala 243:38]
  wire  _GEN_1205 = 3'h5 == io_rob_allocate_allocate_info_bits_1_rob_idx ? 1'h0 : _GEN_1037; // @[Rob.scala 243:38 Rob.scala 243:38]
  wire  _GEN_1206 = 3'h6 == io_rob_allocate_allocate_info_bits_1_rob_idx ? 1'h0 : _GEN_1038; // @[Rob.scala 243:38 Rob.scala 243:38]
  wire  _GEN_1207 = 3'h7 == io_rob_allocate_allocate_info_bits_1_rob_idx ? 1'h0 : _GEN_1039; // @[Rob.scala 243:38 Rob.scala 243:38]
  wire  _GEN_1208 = 3'h0 == io_rob_allocate_allocate_info_bits_1_rob_idx ? 1'h0 : _GEN_1040; // @[Rob.scala 244:30 Rob.scala 244:30]
  wire  _GEN_1209 = 3'h1 == io_rob_allocate_allocate_info_bits_1_rob_idx ? 1'h0 : _GEN_1041; // @[Rob.scala 244:30 Rob.scala 244:30]
  wire  _GEN_1210 = 3'h2 == io_rob_allocate_allocate_info_bits_1_rob_idx ? 1'h0 : _GEN_1042; // @[Rob.scala 244:30 Rob.scala 244:30]
  wire  _GEN_1211 = 3'h3 == io_rob_allocate_allocate_info_bits_1_rob_idx ? 1'h0 : _GEN_1043; // @[Rob.scala 244:30 Rob.scala 244:30]
  wire  _GEN_1212 = 3'h4 == io_rob_allocate_allocate_info_bits_1_rob_idx ? 1'h0 : _GEN_1044; // @[Rob.scala 244:30 Rob.scala 244:30]
  wire  _GEN_1213 = 3'h5 == io_rob_allocate_allocate_info_bits_1_rob_idx ? 1'h0 : _GEN_1045; // @[Rob.scala 244:30 Rob.scala 244:30]
  wire  _GEN_1214 = 3'h6 == io_rob_allocate_allocate_info_bits_1_rob_idx ? 1'h0 : _GEN_1046; // @[Rob.scala 244:30 Rob.scala 244:30]
  wire  _GEN_1215 = 3'h7 == io_rob_allocate_allocate_info_bits_1_rob_idx ? 1'h0 : _GEN_1047; // @[Rob.scala 244:30 Rob.scala 244:30]
  wire  _GEN_1216 = 3'h0 == io_rob_allocate_allocate_info_bits_1_rob_idx | _GEN_1048; // @[Rob.scala 245:34 Rob.scala 245:34]
  wire  _GEN_1217 = 3'h1 == io_rob_allocate_allocate_info_bits_1_rob_idx | _GEN_1049; // @[Rob.scala 245:34 Rob.scala 245:34]
  wire  _GEN_1218 = 3'h2 == io_rob_allocate_allocate_info_bits_1_rob_idx | _GEN_1050; // @[Rob.scala 245:34 Rob.scala 245:34]
  wire  _GEN_1219 = 3'h3 == io_rob_allocate_allocate_info_bits_1_rob_idx | _GEN_1051; // @[Rob.scala 245:34 Rob.scala 245:34]
  wire  _GEN_1220 = 3'h4 == io_rob_allocate_allocate_info_bits_1_rob_idx | _GEN_1052; // @[Rob.scala 245:34 Rob.scala 245:34]
  wire  _GEN_1221 = 3'h5 == io_rob_allocate_allocate_info_bits_1_rob_idx | _GEN_1053; // @[Rob.scala 245:34 Rob.scala 245:34]
  wire  _GEN_1222 = 3'h6 == io_rob_allocate_allocate_info_bits_1_rob_idx | _GEN_1054; // @[Rob.scala 245:34 Rob.scala 245:34]
  wire  _GEN_1223 = 3'h7 == io_rob_allocate_allocate_info_bits_1_rob_idx | _GEN_1055; // @[Rob.scala 245:34 Rob.scala 245:34]
  wire  _GEN_1224 = 3'h0 == io_rob_allocate_allocate_info_bits_1_rob_idx ? 1'h0 : _GEN_1056; // @[Rob.scala 246:35 Rob.scala 246:35]
  wire  _GEN_1225 = 3'h1 == io_rob_allocate_allocate_info_bits_1_rob_idx ? 1'h0 : _GEN_1057; // @[Rob.scala 246:35 Rob.scala 246:35]
  wire  _GEN_1226 = 3'h2 == io_rob_allocate_allocate_info_bits_1_rob_idx ? 1'h0 : _GEN_1058; // @[Rob.scala 246:35 Rob.scala 246:35]
  wire  _GEN_1227 = 3'h3 == io_rob_allocate_allocate_info_bits_1_rob_idx ? 1'h0 : _GEN_1059; // @[Rob.scala 246:35 Rob.scala 246:35]
  wire  _GEN_1228 = 3'h4 == io_rob_allocate_allocate_info_bits_1_rob_idx ? 1'h0 : _GEN_1060; // @[Rob.scala 246:35 Rob.scala 246:35]
  wire  _GEN_1229 = 3'h5 == io_rob_allocate_allocate_info_bits_1_rob_idx ? 1'h0 : _GEN_1061; // @[Rob.scala 246:35 Rob.scala 246:35]
  wire  _GEN_1230 = 3'h6 == io_rob_allocate_allocate_info_bits_1_rob_idx ? 1'h0 : _GEN_1062; // @[Rob.scala 246:35 Rob.scala 246:35]
  wire  _GEN_1231 = 3'h7 == io_rob_allocate_allocate_info_bits_1_rob_idx ? 1'h0 : _GEN_1063; // @[Rob.scala 246:35 Rob.scala 246:35]
  wire  _GEN_1232 = 3'h0 == io_rob_allocate_allocate_info_bits_1_rob_idx ? 1'h0 : _GEN_1064; // @[Rob.scala 247:35 Rob.scala 247:35]
  wire  _GEN_1233 = 3'h1 == io_rob_allocate_allocate_info_bits_1_rob_idx ? 1'h0 : _GEN_1065; // @[Rob.scala 247:35 Rob.scala 247:35]
  wire  _GEN_1234 = 3'h2 == io_rob_allocate_allocate_info_bits_1_rob_idx ? 1'h0 : _GEN_1066; // @[Rob.scala 247:35 Rob.scala 247:35]
  wire  _GEN_1235 = 3'h3 == io_rob_allocate_allocate_info_bits_1_rob_idx ? 1'h0 : _GEN_1067; // @[Rob.scala 247:35 Rob.scala 247:35]
  wire  _GEN_1236 = 3'h4 == io_rob_allocate_allocate_info_bits_1_rob_idx ? 1'h0 : _GEN_1068; // @[Rob.scala 247:35 Rob.scala 247:35]
  wire  _GEN_1237 = 3'h5 == io_rob_allocate_allocate_info_bits_1_rob_idx ? 1'h0 : _GEN_1069; // @[Rob.scala 247:35 Rob.scala 247:35]
  wire  _GEN_1238 = 3'h6 == io_rob_allocate_allocate_info_bits_1_rob_idx ? 1'h0 : _GEN_1070; // @[Rob.scala 247:35 Rob.scala 247:35]
  wire  _GEN_1239 = 3'h7 == io_rob_allocate_allocate_info_bits_1_rob_idx ? 1'h0 : _GEN_1071; // @[Rob.scala 247:35 Rob.scala 247:35]
  wire  _GEN_1240 = 3'h0 == io_rob_allocate_allocate_info_bits_1_rob_idx ? 1'h0 : _GEN_1072; // @[Rob.scala 248:38 Rob.scala 248:38]
  wire  _GEN_1241 = 3'h1 == io_rob_allocate_allocate_info_bits_1_rob_idx ? 1'h0 : _GEN_1073; // @[Rob.scala 248:38 Rob.scala 248:38]
  wire  _GEN_1242 = 3'h2 == io_rob_allocate_allocate_info_bits_1_rob_idx ? 1'h0 : _GEN_1074; // @[Rob.scala 248:38 Rob.scala 248:38]
  wire  _GEN_1243 = 3'h3 == io_rob_allocate_allocate_info_bits_1_rob_idx ? 1'h0 : _GEN_1075; // @[Rob.scala 248:38 Rob.scala 248:38]
  wire  _GEN_1244 = 3'h4 == io_rob_allocate_allocate_info_bits_1_rob_idx ? 1'h0 : _GEN_1076; // @[Rob.scala 248:38 Rob.scala 248:38]
  wire  _GEN_1245 = 3'h5 == io_rob_allocate_allocate_info_bits_1_rob_idx ? 1'h0 : _GEN_1077; // @[Rob.scala 248:38 Rob.scala 248:38]
  wire  _GEN_1246 = 3'h6 == io_rob_allocate_allocate_info_bits_1_rob_idx ? 1'h0 : _GEN_1078; // @[Rob.scala 248:38 Rob.scala 248:38]
  wire  _GEN_1247 = 3'h7 == io_rob_allocate_allocate_info_bits_1_rob_idx ? 1'h0 : _GEN_1079; // @[Rob.scala 248:38 Rob.scala 248:38]
  wire  _GEN_1248 = 3'h0 == io_rob_allocate_allocate_info_bits_1_rob_idx ? 1'h0 : _GEN_1080; // @[Rob.scala 249:34 Rob.scala 249:34]
  wire  _GEN_1249 = 3'h1 == io_rob_allocate_allocate_info_bits_1_rob_idx ? 1'h0 : _GEN_1081; // @[Rob.scala 249:34 Rob.scala 249:34]
  wire  _GEN_1250 = 3'h2 == io_rob_allocate_allocate_info_bits_1_rob_idx ? 1'h0 : _GEN_1082; // @[Rob.scala 249:34 Rob.scala 249:34]
  wire  _GEN_1251 = 3'h3 == io_rob_allocate_allocate_info_bits_1_rob_idx ? 1'h0 : _GEN_1083; // @[Rob.scala 249:34 Rob.scala 249:34]
  wire  _GEN_1252 = 3'h4 == io_rob_allocate_allocate_info_bits_1_rob_idx ? 1'h0 : _GEN_1084; // @[Rob.scala 249:34 Rob.scala 249:34]
  wire  _GEN_1253 = 3'h5 == io_rob_allocate_allocate_info_bits_1_rob_idx ? 1'h0 : _GEN_1085; // @[Rob.scala 249:34 Rob.scala 249:34]
  wire  _GEN_1254 = 3'h6 == io_rob_allocate_allocate_info_bits_1_rob_idx ? 1'h0 : _GEN_1086; // @[Rob.scala 249:34 Rob.scala 249:34]
  wire  _GEN_1255 = 3'h7 == io_rob_allocate_allocate_info_bits_1_rob_idx ? 1'h0 : _GEN_1087; // @[Rob.scala 249:34 Rob.scala 249:34]
  wire  _GEN_1256 = 3'h0 == io_rob_allocate_allocate_info_bits_1_rob_idx ? 1'h0 : _GEN_1088; // @[Rob.scala 250:33 Rob.scala 250:33]
  wire  _GEN_1257 = 3'h1 == io_rob_allocate_allocate_info_bits_1_rob_idx ? 1'h0 : _GEN_1089; // @[Rob.scala 250:33 Rob.scala 250:33]
  wire  _GEN_1258 = 3'h2 == io_rob_allocate_allocate_info_bits_1_rob_idx ? 1'h0 : _GEN_1090; // @[Rob.scala 250:33 Rob.scala 250:33]
  wire  _GEN_1259 = 3'h3 == io_rob_allocate_allocate_info_bits_1_rob_idx ? 1'h0 : _GEN_1091; // @[Rob.scala 250:33 Rob.scala 250:33]
  wire  _GEN_1260 = 3'h4 == io_rob_allocate_allocate_info_bits_1_rob_idx ? 1'h0 : _GEN_1092; // @[Rob.scala 250:33 Rob.scala 250:33]
  wire  _GEN_1261 = 3'h5 == io_rob_allocate_allocate_info_bits_1_rob_idx ? 1'h0 : _GEN_1093; // @[Rob.scala 250:33 Rob.scala 250:33]
  wire  _GEN_1262 = 3'h6 == io_rob_allocate_allocate_info_bits_1_rob_idx ? 1'h0 : _GEN_1094; // @[Rob.scala 250:33 Rob.scala 250:33]
  wire  _GEN_1263 = 3'h7 == io_rob_allocate_allocate_info_bits_1_rob_idx ? 1'h0 : _GEN_1095; // @[Rob.scala 250:33 Rob.scala 250:33]
  wire [31:0] _GEN_1264 = 3'h0 == io_rob_allocate_allocate_info_bits_1_rob_idx ?
    io_rob_allocate_allocate_info_bits_1_inst_addr : _GEN_1096; // @[Rob.scala 251:35 Rob.scala 251:35]
  wire [31:0] _GEN_1265 = 3'h1 == io_rob_allocate_allocate_info_bits_1_rob_idx ?
    io_rob_allocate_allocate_info_bits_1_inst_addr : _GEN_1097; // @[Rob.scala 251:35 Rob.scala 251:35]
  wire [31:0] _GEN_1266 = 3'h2 == io_rob_allocate_allocate_info_bits_1_rob_idx ?
    io_rob_allocate_allocate_info_bits_1_inst_addr : _GEN_1098; // @[Rob.scala 251:35 Rob.scala 251:35]
  wire [31:0] _GEN_1267 = 3'h3 == io_rob_allocate_allocate_info_bits_1_rob_idx ?
    io_rob_allocate_allocate_info_bits_1_inst_addr : _GEN_1099; // @[Rob.scala 251:35 Rob.scala 251:35]
  wire [31:0] _GEN_1268 = 3'h4 == io_rob_allocate_allocate_info_bits_1_rob_idx ?
    io_rob_allocate_allocate_info_bits_1_inst_addr : _GEN_1100; // @[Rob.scala 251:35 Rob.scala 251:35]
  wire [31:0] _GEN_1269 = 3'h5 == io_rob_allocate_allocate_info_bits_1_rob_idx ?
    io_rob_allocate_allocate_info_bits_1_inst_addr : _GEN_1101; // @[Rob.scala 251:35 Rob.scala 251:35]
  wire [31:0] _GEN_1270 = 3'h6 == io_rob_allocate_allocate_info_bits_1_rob_idx ?
    io_rob_allocate_allocate_info_bits_1_inst_addr : _GEN_1102; // @[Rob.scala 251:35 Rob.scala 251:35]
  wire [31:0] _GEN_1271 = 3'h7 == io_rob_allocate_allocate_info_bits_1_rob_idx ?
    io_rob_allocate_allocate_info_bits_1_inst_addr : _GEN_1103; // @[Rob.scala 251:35 Rob.scala 251:35]
  wire [4:0] _GEN_1272 = 3'h0 == io_rob_allocate_allocate_info_bits_1_rob_idx ?
    io_rob_allocate_allocate_info_bits_1_commit_addr[4:0] : _GEN_1104; // @[Rob.scala 252:37 Rob.scala 252:37]
  wire [4:0] _GEN_1273 = 3'h1 == io_rob_allocate_allocate_info_bits_1_rob_idx ?
    io_rob_allocate_allocate_info_bits_1_commit_addr[4:0] : _GEN_1105; // @[Rob.scala 252:37 Rob.scala 252:37]
  wire [4:0] _GEN_1274 = 3'h2 == io_rob_allocate_allocate_info_bits_1_rob_idx ?
    io_rob_allocate_allocate_info_bits_1_commit_addr[4:0] : _GEN_1106; // @[Rob.scala 252:37 Rob.scala 252:37]
  wire [4:0] _GEN_1275 = 3'h3 == io_rob_allocate_allocate_info_bits_1_rob_idx ?
    io_rob_allocate_allocate_info_bits_1_commit_addr[4:0] : _GEN_1107; // @[Rob.scala 252:37 Rob.scala 252:37]
  wire [4:0] _GEN_1276 = 3'h4 == io_rob_allocate_allocate_info_bits_1_rob_idx ?
    io_rob_allocate_allocate_info_bits_1_commit_addr[4:0] : _GEN_1108; // @[Rob.scala 252:37 Rob.scala 252:37]
  wire [4:0] _GEN_1277 = 3'h5 == io_rob_allocate_allocate_info_bits_1_rob_idx ?
    io_rob_allocate_allocate_info_bits_1_commit_addr[4:0] : _GEN_1109; // @[Rob.scala 252:37 Rob.scala 252:37]
  wire [4:0] _GEN_1278 = 3'h6 == io_rob_allocate_allocate_info_bits_1_rob_idx ?
    io_rob_allocate_allocate_info_bits_1_commit_addr[4:0] : _GEN_1110; // @[Rob.scala 252:37 Rob.scala 252:37]
  wire [4:0] _GEN_1279 = 3'h7 == io_rob_allocate_allocate_info_bits_1_rob_idx ?
    io_rob_allocate_allocate_info_bits_1_commit_addr[4:0] : _GEN_1111; // @[Rob.scala 252:37 Rob.scala 252:37]
  wire  _GEN_1296 = 3'h0 == io_rob_allocate_allocate_info_bits_1_rob_idx ? io_rob_allocate_allocate_info_bits_1_unit_sel
     == 3'h5 : _GEN_1128; // @[Rob.scala 255:35 Rob.scala 255:35]
  wire  _GEN_1297 = 3'h1 == io_rob_allocate_allocate_info_bits_1_rob_idx ? io_rob_allocate_allocate_info_bits_1_unit_sel
     == 3'h5 : _GEN_1129; // @[Rob.scala 255:35 Rob.scala 255:35]
  wire  _GEN_1298 = 3'h2 == io_rob_allocate_allocate_info_bits_1_rob_idx ? io_rob_allocate_allocate_info_bits_1_unit_sel
     == 3'h5 : _GEN_1130; // @[Rob.scala 255:35 Rob.scala 255:35]
  wire  _GEN_1299 = 3'h3 == io_rob_allocate_allocate_info_bits_1_rob_idx ? io_rob_allocate_allocate_info_bits_1_unit_sel
     == 3'h5 : _GEN_1131; // @[Rob.scala 255:35 Rob.scala 255:35]
  wire  _GEN_1300 = 3'h4 == io_rob_allocate_allocate_info_bits_1_rob_idx ? io_rob_allocate_allocate_info_bits_1_unit_sel
     == 3'h5 : _GEN_1132; // @[Rob.scala 255:35 Rob.scala 255:35]
  wire  _GEN_1301 = 3'h5 == io_rob_allocate_allocate_info_bits_1_rob_idx ? io_rob_allocate_allocate_info_bits_1_unit_sel
     == 3'h5 : _GEN_1133; // @[Rob.scala 255:35 Rob.scala 255:35]
  wire  _GEN_1302 = 3'h6 == io_rob_allocate_allocate_info_bits_1_rob_idx ? io_rob_allocate_allocate_info_bits_1_unit_sel
     == 3'h5 : _GEN_1134; // @[Rob.scala 255:35 Rob.scala 255:35]
  wire  _GEN_1303 = 3'h7 == io_rob_allocate_allocate_info_bits_1_rob_idx ? io_rob_allocate_allocate_info_bits_1_unit_sel
     == 3'h5 : _GEN_1135; // @[Rob.scala 255:35 Rob.scala 255:35]
  wire [3:0] _GEN_1312 = 3'h0 == io_rob_allocate_allocate_info_bits_1_rob_idx ?
    io_rob_allocate_allocate_info_bits_1_gh_info : _GEN_1144; // @[Rob.scala 257:33 Rob.scala 257:33]
  wire [3:0] _GEN_1313 = 3'h1 == io_rob_allocate_allocate_info_bits_1_rob_idx ?
    io_rob_allocate_allocate_info_bits_1_gh_info : _GEN_1145; // @[Rob.scala 257:33 Rob.scala 257:33]
  wire [3:0] _GEN_1314 = 3'h2 == io_rob_allocate_allocate_info_bits_1_rob_idx ?
    io_rob_allocate_allocate_info_bits_1_gh_info : _GEN_1146; // @[Rob.scala 257:33 Rob.scala 257:33]
  wire [3:0] _GEN_1315 = 3'h3 == io_rob_allocate_allocate_info_bits_1_rob_idx ?
    io_rob_allocate_allocate_info_bits_1_gh_info : _GEN_1147; // @[Rob.scala 257:33 Rob.scala 257:33]
  wire [3:0] _GEN_1316 = 3'h4 == io_rob_allocate_allocate_info_bits_1_rob_idx ?
    io_rob_allocate_allocate_info_bits_1_gh_info : _GEN_1148; // @[Rob.scala 257:33 Rob.scala 257:33]
  wire [3:0] _GEN_1317 = 3'h5 == io_rob_allocate_allocate_info_bits_1_rob_idx ?
    io_rob_allocate_allocate_info_bits_1_gh_info : _GEN_1149; // @[Rob.scala 257:33 Rob.scala 257:33]
  wire [3:0] _GEN_1318 = 3'h6 == io_rob_allocate_allocate_info_bits_1_rob_idx ?
    io_rob_allocate_allocate_info_bits_1_gh_info : _GEN_1150; // @[Rob.scala 257:33 Rob.scala 257:33]
  wire [3:0] _GEN_1319 = 3'h7 == io_rob_allocate_allocate_info_bits_1_rob_idx ?
    io_rob_allocate_allocate_info_bits_1_gh_info : _GEN_1151; // @[Rob.scala 257:33 Rob.scala 257:33]
  wire [5:0] _GEN_1320 = 3'h0 == io_rob_allocate_allocate_info_bits_1_rob_idx ? io_rob_allocate_allocate_info_bits_1_uop
     : _GEN_1152; // @[Rob.scala 258:29 Rob.scala 258:29]
  wire [5:0] _GEN_1321 = 3'h1 == io_rob_allocate_allocate_info_bits_1_rob_idx ? io_rob_allocate_allocate_info_bits_1_uop
     : _GEN_1153; // @[Rob.scala 258:29 Rob.scala 258:29]
  wire [5:0] _GEN_1322 = 3'h2 == io_rob_allocate_allocate_info_bits_1_rob_idx ? io_rob_allocate_allocate_info_bits_1_uop
     : _GEN_1154; // @[Rob.scala 258:29 Rob.scala 258:29]
  wire [5:0] _GEN_1323 = 3'h3 == io_rob_allocate_allocate_info_bits_1_rob_idx ? io_rob_allocate_allocate_info_bits_1_uop
     : _GEN_1155; // @[Rob.scala 258:29 Rob.scala 258:29]
  wire [5:0] _GEN_1324 = 3'h4 == io_rob_allocate_allocate_info_bits_1_rob_idx ? io_rob_allocate_allocate_info_bits_1_uop
     : _GEN_1156; // @[Rob.scala 258:29 Rob.scala 258:29]
  wire [5:0] _GEN_1325 = 3'h5 == io_rob_allocate_allocate_info_bits_1_rob_idx ? io_rob_allocate_allocate_info_bits_1_uop
     : _GEN_1157; // @[Rob.scala 258:29 Rob.scala 258:29]
  wire [5:0] _GEN_1326 = 3'h6 == io_rob_allocate_allocate_info_bits_1_rob_idx ? io_rob_allocate_allocate_info_bits_1_uop
     : _GEN_1158; // @[Rob.scala 258:29 Rob.scala 258:29]
  wire [5:0] _GEN_1327 = 3'h7 == io_rob_allocate_allocate_info_bits_1_rob_idx ? io_rob_allocate_allocate_info_bits_1_uop
     : _GEN_1159; // @[Rob.scala 258:29 Rob.scala 258:29]
  wire [2:0] _GEN_1328 = 3'h0 == io_rob_allocate_allocate_info_bits_1_rob_idx ?
    io_rob_allocate_allocate_info_bits_1_unit_sel : _GEN_1160; // @[Rob.scala 259:34 Rob.scala 259:34]
  wire [2:0] _GEN_1329 = 3'h1 == io_rob_allocate_allocate_info_bits_1_rob_idx ?
    io_rob_allocate_allocate_info_bits_1_unit_sel : _GEN_1161; // @[Rob.scala 259:34 Rob.scala 259:34]
  wire [2:0] _GEN_1330 = 3'h2 == io_rob_allocate_allocate_info_bits_1_rob_idx ?
    io_rob_allocate_allocate_info_bits_1_unit_sel : _GEN_1162; // @[Rob.scala 259:34 Rob.scala 259:34]
  wire [2:0] _GEN_1331 = 3'h3 == io_rob_allocate_allocate_info_bits_1_rob_idx ?
    io_rob_allocate_allocate_info_bits_1_unit_sel : _GEN_1163; // @[Rob.scala 259:34 Rob.scala 259:34]
  wire [2:0] _GEN_1332 = 3'h4 == io_rob_allocate_allocate_info_bits_1_rob_idx ?
    io_rob_allocate_allocate_info_bits_1_unit_sel : _GEN_1164; // @[Rob.scala 259:34 Rob.scala 259:34]
  wire [2:0] _GEN_1333 = 3'h5 == io_rob_allocate_allocate_info_bits_1_rob_idx ?
    io_rob_allocate_allocate_info_bits_1_unit_sel : _GEN_1165; // @[Rob.scala 259:34 Rob.scala 259:34]
  wire [2:0] _GEN_1334 = 3'h6 == io_rob_allocate_allocate_info_bits_1_rob_idx ?
    io_rob_allocate_allocate_info_bits_1_unit_sel : _GEN_1166; // @[Rob.scala 259:34 Rob.scala 259:34]
  wire [2:0] _GEN_1335 = 3'h7 == io_rob_allocate_allocate_info_bits_1_rob_idx ?
    io_rob_allocate_allocate_info_bits_1_unit_sel : _GEN_1167; // @[Rob.scala 259:34 Rob.scala 259:34]
  wire  _GEN_1336 = 3'h0 == io_rob_allocate_allocate_info_bits_1_rob_idx ? io_rob_allocate_allocate_info_bits_1_need_imm
     : _GEN_1168; // @[Rob.scala 260:34 Rob.scala 260:34]
  wire  _GEN_1337 = 3'h1 == io_rob_allocate_allocate_info_bits_1_rob_idx ? io_rob_allocate_allocate_info_bits_1_need_imm
     : _GEN_1169; // @[Rob.scala 260:34 Rob.scala 260:34]
  wire  _GEN_1338 = 3'h2 == io_rob_allocate_allocate_info_bits_1_rob_idx ? io_rob_allocate_allocate_info_bits_1_need_imm
     : _GEN_1170; // @[Rob.scala 260:34 Rob.scala 260:34]
  wire  _GEN_1339 = 3'h3 == io_rob_allocate_allocate_info_bits_1_rob_idx ? io_rob_allocate_allocate_info_bits_1_need_imm
     : _GEN_1171; // @[Rob.scala 260:34 Rob.scala 260:34]
  wire  _GEN_1340 = 3'h4 == io_rob_allocate_allocate_info_bits_1_rob_idx ? io_rob_allocate_allocate_info_bits_1_need_imm
     : _GEN_1172; // @[Rob.scala 260:34 Rob.scala 260:34]
  wire  _GEN_1341 = 3'h5 == io_rob_allocate_allocate_info_bits_1_rob_idx ? io_rob_allocate_allocate_info_bits_1_need_imm
     : _GEN_1173; // @[Rob.scala 260:34 Rob.scala 260:34]
  wire  _GEN_1342 = 3'h6 == io_rob_allocate_allocate_info_bits_1_rob_idx ? io_rob_allocate_allocate_info_bits_1_need_imm
     : _GEN_1174; // @[Rob.scala 260:34 Rob.scala 260:34]
  wire  _GEN_1343 = 3'h7 == io_rob_allocate_allocate_info_bits_1_rob_idx ? io_rob_allocate_allocate_info_bits_1_need_imm
     : _GEN_1175; // @[Rob.scala 260:34 Rob.scala 260:34]
  wire [31:0] _GEN_1344 = 3'h0 == io_rob_allocate_allocate_info_bits_1_rob_idx ?
    io_rob_allocate_allocate_info_bits_1_imm_data : _GEN_1176; // @[Rob.scala 261:34 Rob.scala 261:34]
  wire [31:0] _GEN_1345 = 3'h1 == io_rob_allocate_allocate_info_bits_1_rob_idx ?
    io_rob_allocate_allocate_info_bits_1_imm_data : _GEN_1177; // @[Rob.scala 261:34 Rob.scala 261:34]
  wire [31:0] _GEN_1346 = 3'h2 == io_rob_allocate_allocate_info_bits_1_rob_idx ?
    io_rob_allocate_allocate_info_bits_1_imm_data : _GEN_1178; // @[Rob.scala 261:34 Rob.scala 261:34]
  wire [31:0] _GEN_1347 = 3'h3 == io_rob_allocate_allocate_info_bits_1_rob_idx ?
    io_rob_allocate_allocate_info_bits_1_imm_data : _GEN_1179; // @[Rob.scala 261:34 Rob.scala 261:34]
  wire [31:0] _GEN_1348 = 3'h4 == io_rob_allocate_allocate_info_bits_1_rob_idx ?
    io_rob_allocate_allocate_info_bits_1_imm_data : _GEN_1180; // @[Rob.scala 261:34 Rob.scala 261:34]
  wire [31:0] _GEN_1349 = 3'h5 == io_rob_allocate_allocate_info_bits_1_rob_idx ?
    io_rob_allocate_allocate_info_bits_1_imm_data : _GEN_1181; // @[Rob.scala 261:34 Rob.scala 261:34]
  wire [31:0] _GEN_1350 = 3'h6 == io_rob_allocate_allocate_info_bits_1_rob_idx ?
    io_rob_allocate_allocate_info_bits_1_imm_data : _GEN_1182; // @[Rob.scala 261:34 Rob.scala 261:34]
  wire [31:0] _GEN_1351 = 3'h7 == io_rob_allocate_allocate_info_bits_1_rob_idx ?
    io_rob_allocate_allocate_info_bits_1_imm_data : _GEN_1183; // @[Rob.scala 261:34 Rob.scala 261:34]
  wire  _GEN_1352 = 3'h0 == io_rob_allocate_allocate_info_bits_1_rob_idx ?
    io_rob_allocate_allocate_info_bits_1_flush_on_commit : _GEN_1184; // @[Rob.scala 262:41 Rob.scala 262:41]
  wire  _GEN_1353 = 3'h1 == io_rob_allocate_allocate_info_bits_1_rob_idx ?
    io_rob_allocate_allocate_info_bits_1_flush_on_commit : _GEN_1185; // @[Rob.scala 262:41 Rob.scala 262:41]
  wire  _GEN_1354 = 3'h2 == io_rob_allocate_allocate_info_bits_1_rob_idx ?
    io_rob_allocate_allocate_info_bits_1_flush_on_commit : _GEN_1186; // @[Rob.scala 262:41 Rob.scala 262:41]
  wire  _GEN_1355 = 3'h3 == io_rob_allocate_allocate_info_bits_1_rob_idx ?
    io_rob_allocate_allocate_info_bits_1_flush_on_commit : _GEN_1187; // @[Rob.scala 262:41 Rob.scala 262:41]
  wire  _GEN_1356 = 3'h4 == io_rob_allocate_allocate_info_bits_1_rob_idx ?
    io_rob_allocate_allocate_info_bits_1_flush_on_commit : _GEN_1188; // @[Rob.scala 262:41 Rob.scala 262:41]
  wire  _GEN_1357 = 3'h5 == io_rob_allocate_allocate_info_bits_1_rob_idx ?
    io_rob_allocate_allocate_info_bits_1_flush_on_commit : _GEN_1189; // @[Rob.scala 262:41 Rob.scala 262:41]
  wire  _GEN_1358 = 3'h6 == io_rob_allocate_allocate_info_bits_1_rob_idx ?
    io_rob_allocate_allocate_info_bits_1_flush_on_commit : _GEN_1190; // @[Rob.scala 262:41 Rob.scala 262:41]
  wire  _GEN_1359 = 3'h7 == io_rob_allocate_allocate_info_bits_1_rob_idx ?
    io_rob_allocate_allocate_info_bits_1_flush_on_commit : _GEN_1191; // @[Rob.scala 262:41 Rob.scala 262:41]
  wire  _GEN_1360 = 3'h0 == io_rob_allocate_allocate_info_bits_1_rob_idx ?
    io_rob_allocate_allocate_info_bits_1_predict_taken : _GEN_1192; // @[Rob.scala 263:39 Rob.scala 263:39]
  wire  _GEN_1361 = 3'h1 == io_rob_allocate_allocate_info_bits_1_rob_idx ?
    io_rob_allocate_allocate_info_bits_1_predict_taken : _GEN_1193; // @[Rob.scala 263:39 Rob.scala 263:39]
  wire  _GEN_1362 = 3'h2 == io_rob_allocate_allocate_info_bits_1_rob_idx ?
    io_rob_allocate_allocate_info_bits_1_predict_taken : _GEN_1194; // @[Rob.scala 263:39 Rob.scala 263:39]
  wire  _GEN_1363 = 3'h3 == io_rob_allocate_allocate_info_bits_1_rob_idx ?
    io_rob_allocate_allocate_info_bits_1_predict_taken : _GEN_1195; // @[Rob.scala 263:39 Rob.scala 263:39]
  wire  _GEN_1364 = 3'h4 == io_rob_allocate_allocate_info_bits_1_rob_idx ?
    io_rob_allocate_allocate_info_bits_1_predict_taken : _GEN_1196; // @[Rob.scala 263:39 Rob.scala 263:39]
  wire  _GEN_1365 = 3'h5 == io_rob_allocate_allocate_info_bits_1_rob_idx ?
    io_rob_allocate_allocate_info_bits_1_predict_taken : _GEN_1197; // @[Rob.scala 263:39 Rob.scala 263:39]
  wire  _GEN_1366 = 3'h6 == io_rob_allocate_allocate_info_bits_1_rob_idx ?
    io_rob_allocate_allocate_info_bits_1_predict_taken : _GEN_1198; // @[Rob.scala 263:39 Rob.scala 263:39]
  wire  _GEN_1367 = 3'h7 == io_rob_allocate_allocate_info_bits_1_rob_idx ?
    io_rob_allocate_allocate_info_bits_1_predict_taken : _GEN_1199; // @[Rob.scala 263:39 Rob.scala 263:39]
  wire  _GEN_1368 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1200 : _GEN_1032; // @[Rob.scala 242:112]
  wire  _GEN_1369 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1201 : _GEN_1033; // @[Rob.scala 242:112]
  wire  _GEN_1370 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1202 : _GEN_1034; // @[Rob.scala 242:112]
  wire  _GEN_1371 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1203 : _GEN_1035; // @[Rob.scala 242:112]
  wire  _GEN_1372 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1204 : _GEN_1036; // @[Rob.scala 242:112]
  wire  _GEN_1373 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1205 : _GEN_1037; // @[Rob.scala 242:112]
  wire  _GEN_1374 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1206 : _GEN_1038; // @[Rob.scala 242:112]
  wire  _GEN_1375 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1207 : _GEN_1039; // @[Rob.scala 242:112]
  wire  _GEN_1376 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1208 : _GEN_1040; // @[Rob.scala 242:112]
  wire  _GEN_1377 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1209 : _GEN_1041; // @[Rob.scala 242:112]
  wire  _GEN_1378 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1210 : _GEN_1042; // @[Rob.scala 242:112]
  wire  _GEN_1379 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1211 : _GEN_1043; // @[Rob.scala 242:112]
  wire  _GEN_1380 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1212 : _GEN_1044; // @[Rob.scala 242:112]
  wire  _GEN_1381 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1213 : _GEN_1045; // @[Rob.scala 242:112]
  wire  _GEN_1382 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1214 : _GEN_1046; // @[Rob.scala 242:112]
  wire  _GEN_1383 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1215 : _GEN_1047; // @[Rob.scala 242:112]
  wire  _GEN_1384 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1216 : _GEN_1048; // @[Rob.scala 242:112]
  wire  _GEN_1385 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1217 : _GEN_1049; // @[Rob.scala 242:112]
  wire  _GEN_1386 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1218 : _GEN_1050; // @[Rob.scala 242:112]
  wire  _GEN_1387 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1219 : _GEN_1051; // @[Rob.scala 242:112]
  wire  _GEN_1388 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1220 : _GEN_1052; // @[Rob.scala 242:112]
  wire  _GEN_1389 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1221 : _GEN_1053; // @[Rob.scala 242:112]
  wire  _GEN_1390 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1222 : _GEN_1054; // @[Rob.scala 242:112]
  wire  _GEN_1391 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1223 : _GEN_1055; // @[Rob.scala 242:112]
  wire  _GEN_1392 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1224 : _GEN_1056; // @[Rob.scala 242:112]
  wire  _GEN_1393 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1225 : _GEN_1057; // @[Rob.scala 242:112]
  wire  _GEN_1394 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1226 : _GEN_1058; // @[Rob.scala 242:112]
  wire  _GEN_1395 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1227 : _GEN_1059; // @[Rob.scala 242:112]
  wire  _GEN_1396 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1228 : _GEN_1060; // @[Rob.scala 242:112]
  wire  _GEN_1397 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1229 : _GEN_1061; // @[Rob.scala 242:112]
  wire  _GEN_1398 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1230 : _GEN_1062; // @[Rob.scala 242:112]
  wire  _GEN_1399 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1231 : _GEN_1063; // @[Rob.scala 242:112]
  wire  _GEN_1400 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1232 : _GEN_1064; // @[Rob.scala 242:112]
  wire  _GEN_1401 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1233 : _GEN_1065; // @[Rob.scala 242:112]
  wire  _GEN_1402 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1234 : _GEN_1066; // @[Rob.scala 242:112]
  wire  _GEN_1403 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1235 : _GEN_1067; // @[Rob.scala 242:112]
  wire  _GEN_1404 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1236 : _GEN_1068; // @[Rob.scala 242:112]
  wire  _GEN_1405 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1237 : _GEN_1069; // @[Rob.scala 242:112]
  wire  _GEN_1406 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1238 : _GEN_1070; // @[Rob.scala 242:112]
  wire  _GEN_1407 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1239 : _GEN_1071; // @[Rob.scala 242:112]
  wire  _GEN_1408 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1240 : _GEN_1072; // @[Rob.scala 242:112]
  wire  _GEN_1409 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1241 : _GEN_1073; // @[Rob.scala 242:112]
  wire  _GEN_1410 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1242 : _GEN_1074; // @[Rob.scala 242:112]
  wire  _GEN_1411 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1243 : _GEN_1075; // @[Rob.scala 242:112]
  wire  _GEN_1412 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1244 : _GEN_1076; // @[Rob.scala 242:112]
  wire  _GEN_1413 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1245 : _GEN_1077; // @[Rob.scala 242:112]
  wire  _GEN_1414 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1246 : _GEN_1078; // @[Rob.scala 242:112]
  wire  _GEN_1415 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1247 : _GEN_1079; // @[Rob.scala 242:112]
  wire  _GEN_1416 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1248 : _GEN_1080; // @[Rob.scala 242:112]
  wire  _GEN_1417 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1249 : _GEN_1081; // @[Rob.scala 242:112]
  wire  _GEN_1418 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1250 : _GEN_1082; // @[Rob.scala 242:112]
  wire  _GEN_1419 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1251 : _GEN_1083; // @[Rob.scala 242:112]
  wire  _GEN_1420 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1252 : _GEN_1084; // @[Rob.scala 242:112]
  wire  _GEN_1421 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1253 : _GEN_1085; // @[Rob.scala 242:112]
  wire  _GEN_1422 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1254 : _GEN_1086; // @[Rob.scala 242:112]
  wire  _GEN_1423 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1255 : _GEN_1087; // @[Rob.scala 242:112]
  wire  _GEN_1424 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1256 : _GEN_1088; // @[Rob.scala 242:112]
  wire  _GEN_1425 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1257 : _GEN_1089; // @[Rob.scala 242:112]
  wire  _GEN_1426 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1258 : _GEN_1090; // @[Rob.scala 242:112]
  wire  _GEN_1427 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1259 : _GEN_1091; // @[Rob.scala 242:112]
  wire  _GEN_1428 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1260 : _GEN_1092; // @[Rob.scala 242:112]
  wire  _GEN_1429 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1261 : _GEN_1093; // @[Rob.scala 242:112]
  wire  _GEN_1430 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1262 : _GEN_1094; // @[Rob.scala 242:112]
  wire  _GEN_1431 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1263 : _GEN_1095; // @[Rob.scala 242:112]
  wire [31:0] _GEN_1432 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21
     ? _GEN_1264 : _GEN_1096; // @[Rob.scala 242:112]
  wire [31:0] _GEN_1433 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21
     ? _GEN_1265 : _GEN_1097; // @[Rob.scala 242:112]
  wire [31:0] _GEN_1434 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21
     ? _GEN_1266 : _GEN_1098; // @[Rob.scala 242:112]
  wire [31:0] _GEN_1435 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21
     ? _GEN_1267 : _GEN_1099; // @[Rob.scala 242:112]
  wire [31:0] _GEN_1436 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21
     ? _GEN_1268 : _GEN_1100; // @[Rob.scala 242:112]
  wire [31:0] _GEN_1437 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21
     ? _GEN_1269 : _GEN_1101; // @[Rob.scala 242:112]
  wire [31:0] _GEN_1438 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21
     ? _GEN_1270 : _GEN_1102; // @[Rob.scala 242:112]
  wire [31:0] _GEN_1439 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21
     ? _GEN_1271 : _GEN_1103; // @[Rob.scala 242:112]
  wire [4:0] _GEN_1440 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21
     ? _GEN_1272 : _GEN_1104; // @[Rob.scala 242:112]
  wire [4:0] _GEN_1441 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21
     ? _GEN_1273 : _GEN_1105; // @[Rob.scala 242:112]
  wire [4:0] _GEN_1442 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21
     ? _GEN_1274 : _GEN_1106; // @[Rob.scala 242:112]
  wire [4:0] _GEN_1443 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21
     ? _GEN_1275 : _GEN_1107; // @[Rob.scala 242:112]
  wire [4:0] _GEN_1444 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21
     ? _GEN_1276 : _GEN_1108; // @[Rob.scala 242:112]
  wire [4:0] _GEN_1445 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21
     ? _GEN_1277 : _GEN_1109; // @[Rob.scala 242:112]
  wire [4:0] _GEN_1446 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21
     ? _GEN_1278 : _GEN_1110; // @[Rob.scala 242:112]
  wire [4:0] _GEN_1447 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21
     ? _GEN_1279 : _GEN_1111; // @[Rob.scala 242:112]
  wire  _GEN_1464 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1296 : _GEN_1128; // @[Rob.scala 242:112]
  wire  _GEN_1465 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1297 : _GEN_1129; // @[Rob.scala 242:112]
  wire  _GEN_1466 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1298 : _GEN_1130; // @[Rob.scala 242:112]
  wire  _GEN_1467 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1299 : _GEN_1131; // @[Rob.scala 242:112]
  wire  _GEN_1468 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1300 : _GEN_1132; // @[Rob.scala 242:112]
  wire  _GEN_1469 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1301 : _GEN_1133; // @[Rob.scala 242:112]
  wire  _GEN_1470 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1302 : _GEN_1134; // @[Rob.scala 242:112]
  wire  _GEN_1471 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1303 : _GEN_1135; // @[Rob.scala 242:112]
  wire [3:0] _GEN_1480 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21
     ? _GEN_1312 : _GEN_1144; // @[Rob.scala 242:112]
  wire [3:0] _GEN_1481 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21
     ? _GEN_1313 : _GEN_1145; // @[Rob.scala 242:112]
  wire [3:0] _GEN_1482 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21
     ? _GEN_1314 : _GEN_1146; // @[Rob.scala 242:112]
  wire [3:0] _GEN_1483 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21
     ? _GEN_1315 : _GEN_1147; // @[Rob.scala 242:112]
  wire [3:0] _GEN_1484 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21
     ? _GEN_1316 : _GEN_1148; // @[Rob.scala 242:112]
  wire [3:0] _GEN_1485 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21
     ? _GEN_1317 : _GEN_1149; // @[Rob.scala 242:112]
  wire [3:0] _GEN_1486 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21
     ? _GEN_1318 : _GEN_1150; // @[Rob.scala 242:112]
  wire [3:0] _GEN_1487 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21
     ? _GEN_1319 : _GEN_1151; // @[Rob.scala 242:112]
  wire [5:0] _GEN_1488 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21
     ? _GEN_1320 : _GEN_1152; // @[Rob.scala 242:112]
  wire [5:0] _GEN_1489 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21
     ? _GEN_1321 : _GEN_1153; // @[Rob.scala 242:112]
  wire [5:0] _GEN_1490 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21
     ? _GEN_1322 : _GEN_1154; // @[Rob.scala 242:112]
  wire [5:0] _GEN_1491 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21
     ? _GEN_1323 : _GEN_1155; // @[Rob.scala 242:112]
  wire [5:0] _GEN_1492 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21
     ? _GEN_1324 : _GEN_1156; // @[Rob.scala 242:112]
  wire [5:0] _GEN_1493 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21
     ? _GEN_1325 : _GEN_1157; // @[Rob.scala 242:112]
  wire [5:0] _GEN_1494 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21
     ? _GEN_1326 : _GEN_1158; // @[Rob.scala 242:112]
  wire [5:0] _GEN_1495 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21
     ? _GEN_1327 : _GEN_1159; // @[Rob.scala 242:112]
  wire [2:0] _GEN_1496 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21
     ? _GEN_1328 : _GEN_1160; // @[Rob.scala 242:112]
  wire [2:0] _GEN_1497 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21
     ? _GEN_1329 : _GEN_1161; // @[Rob.scala 242:112]
  wire [2:0] _GEN_1498 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21
     ? _GEN_1330 : _GEN_1162; // @[Rob.scala 242:112]
  wire [2:0] _GEN_1499 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21
     ? _GEN_1331 : _GEN_1163; // @[Rob.scala 242:112]
  wire [2:0] _GEN_1500 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21
     ? _GEN_1332 : _GEN_1164; // @[Rob.scala 242:112]
  wire [2:0] _GEN_1501 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21
     ? _GEN_1333 : _GEN_1165; // @[Rob.scala 242:112]
  wire [2:0] _GEN_1502 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21
     ? _GEN_1334 : _GEN_1166; // @[Rob.scala 242:112]
  wire [2:0] _GEN_1503 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21
     ? _GEN_1335 : _GEN_1167; // @[Rob.scala 242:112]
  wire  _GEN_1504 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1336 : _GEN_1168; // @[Rob.scala 242:112]
  wire  _GEN_1505 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1337 : _GEN_1169; // @[Rob.scala 242:112]
  wire  _GEN_1506 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1338 : _GEN_1170; // @[Rob.scala 242:112]
  wire  _GEN_1507 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1339 : _GEN_1171; // @[Rob.scala 242:112]
  wire  _GEN_1508 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1340 : _GEN_1172; // @[Rob.scala 242:112]
  wire  _GEN_1509 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1341 : _GEN_1173; // @[Rob.scala 242:112]
  wire  _GEN_1510 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1342 : _GEN_1174; // @[Rob.scala 242:112]
  wire  _GEN_1511 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1343 : _GEN_1175; // @[Rob.scala 242:112]
  wire [31:0] _GEN_1512 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21
     ? _GEN_1344 : _GEN_1176; // @[Rob.scala 242:112]
  wire [31:0] _GEN_1513 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21
     ? _GEN_1345 : _GEN_1177; // @[Rob.scala 242:112]
  wire [31:0] _GEN_1514 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21
     ? _GEN_1346 : _GEN_1178; // @[Rob.scala 242:112]
  wire [31:0] _GEN_1515 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21
     ? _GEN_1347 : _GEN_1179; // @[Rob.scala 242:112]
  wire [31:0] _GEN_1516 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21
     ? _GEN_1348 : _GEN_1180; // @[Rob.scala 242:112]
  wire [31:0] _GEN_1517 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21
     ? _GEN_1349 : _GEN_1181; // @[Rob.scala 242:112]
  wire [31:0] _GEN_1518 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21
     ? _GEN_1350 : _GEN_1182; // @[Rob.scala 242:112]
  wire [31:0] _GEN_1519 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21
     ? _GEN_1351 : _GEN_1183; // @[Rob.scala 242:112]
  wire  _GEN_1520 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1352 : _GEN_1184; // @[Rob.scala 242:112]
  wire  _GEN_1521 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1353 : _GEN_1185; // @[Rob.scala 242:112]
  wire  _GEN_1522 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1354 : _GEN_1186; // @[Rob.scala 242:112]
  wire  _GEN_1523 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1355 : _GEN_1187; // @[Rob.scala 242:112]
  wire  _GEN_1524 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1356 : _GEN_1188; // @[Rob.scala 242:112]
  wire  _GEN_1525 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1357 : _GEN_1189; // @[Rob.scala 242:112]
  wire  _GEN_1526 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1358 : _GEN_1190; // @[Rob.scala 242:112]
  wire  _GEN_1527 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1359 : _GEN_1191; // @[Rob.scala 242:112]
  wire  _GEN_1528 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1360 : _GEN_1192; // @[Rob.scala 242:112]
  wire  _GEN_1529 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1361 : _GEN_1193; // @[Rob.scala 242:112]
  wire  _GEN_1530 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1362 : _GEN_1194; // @[Rob.scala 242:112]
  wire  _GEN_1531 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1363 : _GEN_1195; // @[Rob.scala 242:112]
  wire  _GEN_1532 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1364 : _GEN_1196; // @[Rob.scala 242:112]
  wire  _GEN_1533 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1365 : _GEN_1197; // @[Rob.scala 242:112]
  wire  _GEN_1534 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1366 : _GEN_1198; // @[Rob.scala 242:112]
  wire  _GEN_1535 = io_rob_allocate_allocate_info_valid & io_rob_allocate_allocate_info_bits_1_inst_valid & _T_21 ?
    _GEN_1367 : _GEN_1199; // @[Rob.scala 242:112]
  wire [31:0] _GEN_1536 = io_wb_info_i_0_valid & io_wb_info_i_0_bits_rob_idx == rob_info_0_op1_tag & rob_info_0_is_valid
     & ~rob_info_0_op1_ready & rob_info_0_is_init & _T_21 ? io_wb_info_i_0_bits_data : rob_info_0_op1_data; // @[Rob.scala 269:177 Rob.scala 270:30 Rob.scala 175:27]
  wire [31:0] _GEN_1538 = io_wb_info_i_0_valid & io_wb_info_i_0_bits_rob_idx == rob_info_0_op2_tag & rob_info_0_is_valid
     & ~rob_info_0_op2_ready & rob_info_0_is_init & _T_21 ? io_wb_info_i_0_bits_data : rob_info_0_op2_data; // @[Rob.scala 273:177 Rob.scala 274:30 Rob.scala 175:27]
  wire [31:0] _GEN_1540 = io_wb_info_i_1_valid & io_wb_info_i_1_bits_rob_idx == rob_info_0_op1_tag & rob_info_0_is_valid
     & ~rob_info_0_op1_ready & rob_info_0_is_init & _T_21 ? io_wb_info_i_1_bits_data : _GEN_1536; // @[Rob.scala 269:177 Rob.scala 270:30]
  wire [31:0] _GEN_1542 = io_wb_info_i_1_valid & io_wb_info_i_1_bits_rob_idx == rob_info_0_op2_tag & rob_info_0_is_valid
     & ~rob_info_0_op2_ready & rob_info_0_is_init & _T_21 ? io_wb_info_i_1_bits_data : _GEN_1538; // @[Rob.scala 273:177 Rob.scala 274:30]
  wire [31:0] _GEN_1544 = io_wb_info_i_2_valid & io_wb_info_i_2_bits_rob_idx == rob_info_0_op1_tag & rob_info_0_is_valid
     & ~rob_info_0_op1_ready & rob_info_0_is_init & _T_21 ? io_wb_info_i_2_bits_data : _GEN_1540; // @[Rob.scala 269:177 Rob.scala 270:30]
  wire  _GEN_1545 = io_wb_info_i_2_valid & io_wb_info_i_2_bits_rob_idx == rob_info_0_op1_tag & rob_info_0_is_valid & ~
    rob_info_0_op1_ready & rob_info_0_is_init & _T_21 | (io_wb_info_i_1_valid & io_wb_info_i_1_bits_rob_idx ==
    rob_info_0_op1_tag & rob_info_0_is_valid & ~rob_info_0_op1_ready & rob_info_0_is_init & _T_21 | (
    io_wb_info_i_0_valid & io_wb_info_i_0_bits_rob_idx == rob_info_0_op1_tag & rob_info_0_is_valid & ~
    rob_info_0_op1_ready & rob_info_0_is_init & _T_21 | _GEN_1392)); // @[Rob.scala 269:177 Rob.scala 271:31]
  wire [31:0] _GEN_1546 = io_wb_info_i_2_valid & io_wb_info_i_2_bits_rob_idx == rob_info_0_op2_tag & rob_info_0_is_valid
     & ~rob_info_0_op2_ready & rob_info_0_is_init & _T_21 ? io_wb_info_i_2_bits_data : _GEN_1542; // @[Rob.scala 273:177 Rob.scala 274:30]
  wire  _GEN_1547 = io_wb_info_i_2_valid & io_wb_info_i_2_bits_rob_idx == rob_info_0_op2_tag & rob_info_0_is_valid & ~
    rob_info_0_op2_ready & rob_info_0_is_init & _T_21 | (io_wb_info_i_1_valid & io_wb_info_i_1_bits_rob_idx ==
    rob_info_0_op2_tag & rob_info_0_is_valid & ~rob_info_0_op2_ready & rob_info_0_is_init & _T_21 | (
    io_wb_info_i_0_valid & io_wb_info_i_0_bits_rob_idx == rob_info_0_op2_tag & rob_info_0_is_valid & ~
    rob_info_0_op2_ready & rob_info_0_is_init & _T_21 | _GEN_1400)); // @[Rob.scala 273:177 Rob.scala 275:31]
  wire [31:0] _GEN_1548 = io_wb_info_i_3_valid & io_wb_info_i_3_bits_rob_idx == rob_info_0_op1_tag & rob_info_0_is_valid
     & ~rob_info_0_op1_ready & rob_info_0_is_init & _T_21 ? io_wb_info_i_3_bits_data : _GEN_1544; // @[Rob.scala 269:177 Rob.scala 270:30]
  wire [31:0] _GEN_1550 = io_wb_info_i_3_valid & io_wb_info_i_3_bits_rob_idx == rob_info_0_op2_tag & rob_info_0_is_valid
     & ~rob_info_0_op2_ready & rob_info_0_is_init & _T_21 ? io_wb_info_i_3_bits_data : _GEN_1546; // @[Rob.scala 273:177 Rob.scala 274:30]
  wire [31:0] _GEN_1552 = io_wb_info_i_4_valid & io_wb_info_i_4_bits_rob_idx == rob_info_0_op1_tag & rob_info_0_is_valid
     & ~rob_info_0_op1_ready & rob_info_0_is_init & _T_21 ? io_wb_info_i_4_bits_data : _GEN_1548; // @[Rob.scala 269:177 Rob.scala 270:30]
  wire  _GEN_1553 = io_wb_info_i_4_valid & io_wb_info_i_4_bits_rob_idx == rob_info_0_op1_tag & rob_info_0_is_valid & ~
    rob_info_0_op1_ready & rob_info_0_is_init & _T_21 | (io_wb_info_i_3_valid & io_wb_info_i_3_bits_rob_idx ==
    rob_info_0_op1_tag & rob_info_0_is_valid & ~rob_info_0_op1_ready & rob_info_0_is_init & _T_21 | _GEN_1545); // @[Rob.scala 269:177 Rob.scala 271:31]
  wire [31:0] _GEN_1554 = io_wb_info_i_4_valid & io_wb_info_i_4_bits_rob_idx == rob_info_0_op2_tag & rob_info_0_is_valid
     & ~rob_info_0_op2_ready & rob_info_0_is_init & _T_21 ? io_wb_info_i_4_bits_data : _GEN_1550; // @[Rob.scala 273:177 Rob.scala 274:30]
  wire  _GEN_1555 = io_wb_info_i_4_valid & io_wb_info_i_4_bits_rob_idx == rob_info_0_op2_tag & rob_info_0_is_valid & ~
    rob_info_0_op2_ready & rob_info_0_is_init & _T_21 | (io_wb_info_i_3_valid & io_wb_info_i_3_bits_rob_idx ==
    rob_info_0_op2_tag & rob_info_0_is_valid & ~rob_info_0_op2_ready & rob_info_0_is_init & _T_21 | _GEN_1547); // @[Rob.scala 273:177 Rob.scala 275:31]
  wire [31:0] _GEN_1556 = io_wb_info_i_0_valid & io_wb_info_i_0_bits_rob_idx == rob_info_1_op1_tag & rob_info_1_is_valid
     & ~rob_info_1_op1_ready & rob_info_1_is_init & _T_21 ? io_wb_info_i_0_bits_data : rob_info_1_op1_data; // @[Rob.scala 269:177 Rob.scala 270:30 Rob.scala 175:27]
  wire [31:0] _GEN_1558 = io_wb_info_i_0_valid & io_wb_info_i_0_bits_rob_idx == rob_info_1_op2_tag & rob_info_1_is_valid
     & ~rob_info_1_op2_ready & rob_info_1_is_init & _T_21 ? io_wb_info_i_0_bits_data : rob_info_1_op2_data; // @[Rob.scala 273:177 Rob.scala 274:30 Rob.scala 175:27]
  wire [31:0] _GEN_1560 = io_wb_info_i_1_valid & io_wb_info_i_1_bits_rob_idx == rob_info_1_op1_tag & rob_info_1_is_valid
     & ~rob_info_1_op1_ready & rob_info_1_is_init & _T_21 ? io_wb_info_i_1_bits_data : _GEN_1556; // @[Rob.scala 269:177 Rob.scala 270:30]
  wire [31:0] _GEN_1562 = io_wb_info_i_1_valid & io_wb_info_i_1_bits_rob_idx == rob_info_1_op2_tag & rob_info_1_is_valid
     & ~rob_info_1_op2_ready & rob_info_1_is_init & _T_21 ? io_wb_info_i_1_bits_data : _GEN_1558; // @[Rob.scala 273:177 Rob.scala 274:30]
  wire [31:0] _GEN_1564 = io_wb_info_i_2_valid & io_wb_info_i_2_bits_rob_idx == rob_info_1_op1_tag & rob_info_1_is_valid
     & ~rob_info_1_op1_ready & rob_info_1_is_init & _T_21 ? io_wb_info_i_2_bits_data : _GEN_1560; // @[Rob.scala 269:177 Rob.scala 270:30]
  wire  _GEN_1565 = io_wb_info_i_2_valid & io_wb_info_i_2_bits_rob_idx == rob_info_1_op1_tag & rob_info_1_is_valid & ~
    rob_info_1_op1_ready & rob_info_1_is_init & _T_21 | (io_wb_info_i_1_valid & io_wb_info_i_1_bits_rob_idx ==
    rob_info_1_op1_tag & rob_info_1_is_valid & ~rob_info_1_op1_ready & rob_info_1_is_init & _T_21 | (
    io_wb_info_i_0_valid & io_wb_info_i_0_bits_rob_idx == rob_info_1_op1_tag & rob_info_1_is_valid & ~
    rob_info_1_op1_ready & rob_info_1_is_init & _T_21 | _GEN_1393)); // @[Rob.scala 269:177 Rob.scala 271:31]
  wire [31:0] _GEN_1566 = io_wb_info_i_2_valid & io_wb_info_i_2_bits_rob_idx == rob_info_1_op2_tag & rob_info_1_is_valid
     & ~rob_info_1_op2_ready & rob_info_1_is_init & _T_21 ? io_wb_info_i_2_bits_data : _GEN_1562; // @[Rob.scala 273:177 Rob.scala 274:30]
  wire  _GEN_1567 = io_wb_info_i_2_valid & io_wb_info_i_2_bits_rob_idx == rob_info_1_op2_tag & rob_info_1_is_valid & ~
    rob_info_1_op2_ready & rob_info_1_is_init & _T_21 | (io_wb_info_i_1_valid & io_wb_info_i_1_bits_rob_idx ==
    rob_info_1_op2_tag & rob_info_1_is_valid & ~rob_info_1_op2_ready & rob_info_1_is_init & _T_21 | (
    io_wb_info_i_0_valid & io_wb_info_i_0_bits_rob_idx == rob_info_1_op2_tag & rob_info_1_is_valid & ~
    rob_info_1_op2_ready & rob_info_1_is_init & _T_21 | _GEN_1401)); // @[Rob.scala 273:177 Rob.scala 275:31]
  wire [31:0] _GEN_1568 = io_wb_info_i_3_valid & io_wb_info_i_3_bits_rob_idx == rob_info_1_op1_tag & rob_info_1_is_valid
     & ~rob_info_1_op1_ready & rob_info_1_is_init & _T_21 ? io_wb_info_i_3_bits_data : _GEN_1564; // @[Rob.scala 269:177 Rob.scala 270:30]
  wire [31:0] _GEN_1570 = io_wb_info_i_3_valid & io_wb_info_i_3_bits_rob_idx == rob_info_1_op2_tag & rob_info_1_is_valid
     & ~rob_info_1_op2_ready & rob_info_1_is_init & _T_21 ? io_wb_info_i_3_bits_data : _GEN_1566; // @[Rob.scala 273:177 Rob.scala 274:30]
  wire [31:0] _GEN_1572 = io_wb_info_i_4_valid & io_wb_info_i_4_bits_rob_idx == rob_info_1_op1_tag & rob_info_1_is_valid
     & ~rob_info_1_op1_ready & rob_info_1_is_init & _T_21 ? io_wb_info_i_4_bits_data : _GEN_1568; // @[Rob.scala 269:177 Rob.scala 270:30]
  wire  _GEN_1573 = io_wb_info_i_4_valid & io_wb_info_i_4_bits_rob_idx == rob_info_1_op1_tag & rob_info_1_is_valid & ~
    rob_info_1_op1_ready & rob_info_1_is_init & _T_21 | (io_wb_info_i_3_valid & io_wb_info_i_3_bits_rob_idx ==
    rob_info_1_op1_tag & rob_info_1_is_valid & ~rob_info_1_op1_ready & rob_info_1_is_init & _T_21 | _GEN_1565); // @[Rob.scala 269:177 Rob.scala 271:31]
  wire [31:0] _GEN_1574 = io_wb_info_i_4_valid & io_wb_info_i_4_bits_rob_idx == rob_info_1_op2_tag & rob_info_1_is_valid
     & ~rob_info_1_op2_ready & rob_info_1_is_init & _T_21 ? io_wb_info_i_4_bits_data : _GEN_1570; // @[Rob.scala 273:177 Rob.scala 274:30]
  wire  _GEN_1575 = io_wb_info_i_4_valid & io_wb_info_i_4_bits_rob_idx == rob_info_1_op2_tag & rob_info_1_is_valid & ~
    rob_info_1_op2_ready & rob_info_1_is_init & _T_21 | (io_wb_info_i_3_valid & io_wb_info_i_3_bits_rob_idx ==
    rob_info_1_op2_tag & rob_info_1_is_valid & ~rob_info_1_op2_ready & rob_info_1_is_init & _T_21 | _GEN_1567); // @[Rob.scala 273:177 Rob.scala 275:31]
  wire [31:0] _GEN_1576 = io_wb_info_i_0_valid & io_wb_info_i_0_bits_rob_idx == rob_info_2_op1_tag & rob_info_2_is_valid
     & ~rob_info_2_op1_ready & rob_info_2_is_init & _T_21 ? io_wb_info_i_0_bits_data : rob_info_2_op1_data; // @[Rob.scala 269:177 Rob.scala 270:30 Rob.scala 175:27]
  wire [31:0] _GEN_1578 = io_wb_info_i_0_valid & io_wb_info_i_0_bits_rob_idx == rob_info_2_op2_tag & rob_info_2_is_valid
     & ~rob_info_2_op2_ready & rob_info_2_is_init & _T_21 ? io_wb_info_i_0_bits_data : rob_info_2_op2_data; // @[Rob.scala 273:177 Rob.scala 274:30 Rob.scala 175:27]
  wire [31:0] _GEN_1580 = io_wb_info_i_1_valid & io_wb_info_i_1_bits_rob_idx == rob_info_2_op1_tag & rob_info_2_is_valid
     & ~rob_info_2_op1_ready & rob_info_2_is_init & _T_21 ? io_wb_info_i_1_bits_data : _GEN_1576; // @[Rob.scala 269:177 Rob.scala 270:30]
  wire [31:0] _GEN_1582 = io_wb_info_i_1_valid & io_wb_info_i_1_bits_rob_idx == rob_info_2_op2_tag & rob_info_2_is_valid
     & ~rob_info_2_op2_ready & rob_info_2_is_init & _T_21 ? io_wb_info_i_1_bits_data : _GEN_1578; // @[Rob.scala 273:177 Rob.scala 274:30]
  wire [31:0] _GEN_1584 = io_wb_info_i_2_valid & io_wb_info_i_2_bits_rob_idx == rob_info_2_op1_tag & rob_info_2_is_valid
     & ~rob_info_2_op1_ready & rob_info_2_is_init & _T_21 ? io_wb_info_i_2_bits_data : _GEN_1580; // @[Rob.scala 269:177 Rob.scala 270:30]
  wire  _GEN_1585 = io_wb_info_i_2_valid & io_wb_info_i_2_bits_rob_idx == rob_info_2_op1_tag & rob_info_2_is_valid & ~
    rob_info_2_op1_ready & rob_info_2_is_init & _T_21 | (io_wb_info_i_1_valid & io_wb_info_i_1_bits_rob_idx ==
    rob_info_2_op1_tag & rob_info_2_is_valid & ~rob_info_2_op1_ready & rob_info_2_is_init & _T_21 | (
    io_wb_info_i_0_valid & io_wb_info_i_0_bits_rob_idx == rob_info_2_op1_tag & rob_info_2_is_valid & ~
    rob_info_2_op1_ready & rob_info_2_is_init & _T_21 | _GEN_1394)); // @[Rob.scala 269:177 Rob.scala 271:31]
  wire [31:0] _GEN_1586 = io_wb_info_i_2_valid & io_wb_info_i_2_bits_rob_idx == rob_info_2_op2_tag & rob_info_2_is_valid
     & ~rob_info_2_op2_ready & rob_info_2_is_init & _T_21 ? io_wb_info_i_2_bits_data : _GEN_1582; // @[Rob.scala 273:177 Rob.scala 274:30]
  wire  _GEN_1587 = io_wb_info_i_2_valid & io_wb_info_i_2_bits_rob_idx == rob_info_2_op2_tag & rob_info_2_is_valid & ~
    rob_info_2_op2_ready & rob_info_2_is_init & _T_21 | (io_wb_info_i_1_valid & io_wb_info_i_1_bits_rob_idx ==
    rob_info_2_op2_tag & rob_info_2_is_valid & ~rob_info_2_op2_ready & rob_info_2_is_init & _T_21 | (
    io_wb_info_i_0_valid & io_wb_info_i_0_bits_rob_idx == rob_info_2_op2_tag & rob_info_2_is_valid & ~
    rob_info_2_op2_ready & rob_info_2_is_init & _T_21 | _GEN_1402)); // @[Rob.scala 273:177 Rob.scala 275:31]
  wire [31:0] _GEN_1588 = io_wb_info_i_3_valid & io_wb_info_i_3_bits_rob_idx == rob_info_2_op1_tag & rob_info_2_is_valid
     & ~rob_info_2_op1_ready & rob_info_2_is_init & _T_21 ? io_wb_info_i_3_bits_data : _GEN_1584; // @[Rob.scala 269:177 Rob.scala 270:30]
  wire [31:0] _GEN_1590 = io_wb_info_i_3_valid & io_wb_info_i_3_bits_rob_idx == rob_info_2_op2_tag & rob_info_2_is_valid
     & ~rob_info_2_op2_ready & rob_info_2_is_init & _T_21 ? io_wb_info_i_3_bits_data : _GEN_1586; // @[Rob.scala 273:177 Rob.scala 274:30]
  wire [31:0] _GEN_1592 = io_wb_info_i_4_valid & io_wb_info_i_4_bits_rob_idx == rob_info_2_op1_tag & rob_info_2_is_valid
     & ~rob_info_2_op1_ready & rob_info_2_is_init & _T_21 ? io_wb_info_i_4_bits_data : _GEN_1588; // @[Rob.scala 269:177 Rob.scala 270:30]
  wire  _GEN_1593 = io_wb_info_i_4_valid & io_wb_info_i_4_bits_rob_idx == rob_info_2_op1_tag & rob_info_2_is_valid & ~
    rob_info_2_op1_ready & rob_info_2_is_init & _T_21 | (io_wb_info_i_3_valid & io_wb_info_i_3_bits_rob_idx ==
    rob_info_2_op1_tag & rob_info_2_is_valid & ~rob_info_2_op1_ready & rob_info_2_is_init & _T_21 | _GEN_1585); // @[Rob.scala 269:177 Rob.scala 271:31]
  wire [31:0] _GEN_1594 = io_wb_info_i_4_valid & io_wb_info_i_4_bits_rob_idx == rob_info_2_op2_tag & rob_info_2_is_valid
     & ~rob_info_2_op2_ready & rob_info_2_is_init & _T_21 ? io_wb_info_i_4_bits_data : _GEN_1590; // @[Rob.scala 273:177 Rob.scala 274:30]
  wire  _GEN_1595 = io_wb_info_i_4_valid & io_wb_info_i_4_bits_rob_idx == rob_info_2_op2_tag & rob_info_2_is_valid & ~
    rob_info_2_op2_ready & rob_info_2_is_init & _T_21 | (io_wb_info_i_3_valid & io_wb_info_i_3_bits_rob_idx ==
    rob_info_2_op2_tag & rob_info_2_is_valid & ~rob_info_2_op2_ready & rob_info_2_is_init & _T_21 | _GEN_1587); // @[Rob.scala 273:177 Rob.scala 275:31]
  wire [31:0] _GEN_1596 = io_wb_info_i_0_valid & io_wb_info_i_0_bits_rob_idx == rob_info_3_op1_tag & rob_info_3_is_valid
     & ~rob_info_3_op1_ready & rob_info_3_is_init & _T_21 ? io_wb_info_i_0_bits_data : rob_info_3_op1_data; // @[Rob.scala 269:177 Rob.scala 270:30 Rob.scala 175:27]
  wire [31:0] _GEN_1598 = io_wb_info_i_0_valid & io_wb_info_i_0_bits_rob_idx == rob_info_3_op2_tag & rob_info_3_is_valid
     & ~rob_info_3_op2_ready & rob_info_3_is_init & _T_21 ? io_wb_info_i_0_bits_data : rob_info_3_op2_data; // @[Rob.scala 273:177 Rob.scala 274:30 Rob.scala 175:27]
  wire [31:0] _GEN_1600 = io_wb_info_i_1_valid & io_wb_info_i_1_bits_rob_idx == rob_info_3_op1_tag & rob_info_3_is_valid
     & ~rob_info_3_op1_ready & rob_info_3_is_init & _T_21 ? io_wb_info_i_1_bits_data : _GEN_1596; // @[Rob.scala 269:177 Rob.scala 270:30]
  wire [31:0] _GEN_1602 = io_wb_info_i_1_valid & io_wb_info_i_1_bits_rob_idx == rob_info_3_op2_tag & rob_info_3_is_valid
     & ~rob_info_3_op2_ready & rob_info_3_is_init & _T_21 ? io_wb_info_i_1_bits_data : _GEN_1598; // @[Rob.scala 273:177 Rob.scala 274:30]
  wire [31:0] _GEN_1604 = io_wb_info_i_2_valid & io_wb_info_i_2_bits_rob_idx == rob_info_3_op1_tag & rob_info_3_is_valid
     & ~rob_info_3_op1_ready & rob_info_3_is_init & _T_21 ? io_wb_info_i_2_bits_data : _GEN_1600; // @[Rob.scala 269:177 Rob.scala 270:30]
  wire  _GEN_1605 = io_wb_info_i_2_valid & io_wb_info_i_2_bits_rob_idx == rob_info_3_op1_tag & rob_info_3_is_valid & ~
    rob_info_3_op1_ready & rob_info_3_is_init & _T_21 | (io_wb_info_i_1_valid & io_wb_info_i_1_bits_rob_idx ==
    rob_info_3_op1_tag & rob_info_3_is_valid & ~rob_info_3_op1_ready & rob_info_3_is_init & _T_21 | (
    io_wb_info_i_0_valid & io_wb_info_i_0_bits_rob_idx == rob_info_3_op1_tag & rob_info_3_is_valid & ~
    rob_info_3_op1_ready & rob_info_3_is_init & _T_21 | _GEN_1395)); // @[Rob.scala 269:177 Rob.scala 271:31]
  wire [31:0] _GEN_1606 = io_wb_info_i_2_valid & io_wb_info_i_2_bits_rob_idx == rob_info_3_op2_tag & rob_info_3_is_valid
     & ~rob_info_3_op2_ready & rob_info_3_is_init & _T_21 ? io_wb_info_i_2_bits_data : _GEN_1602; // @[Rob.scala 273:177 Rob.scala 274:30]
  wire  _GEN_1607 = io_wb_info_i_2_valid & io_wb_info_i_2_bits_rob_idx == rob_info_3_op2_tag & rob_info_3_is_valid & ~
    rob_info_3_op2_ready & rob_info_3_is_init & _T_21 | (io_wb_info_i_1_valid & io_wb_info_i_1_bits_rob_idx ==
    rob_info_3_op2_tag & rob_info_3_is_valid & ~rob_info_3_op2_ready & rob_info_3_is_init & _T_21 | (
    io_wb_info_i_0_valid & io_wb_info_i_0_bits_rob_idx == rob_info_3_op2_tag & rob_info_3_is_valid & ~
    rob_info_3_op2_ready & rob_info_3_is_init & _T_21 | _GEN_1403)); // @[Rob.scala 273:177 Rob.scala 275:31]
  wire [31:0] _GEN_1608 = io_wb_info_i_3_valid & io_wb_info_i_3_bits_rob_idx == rob_info_3_op1_tag & rob_info_3_is_valid
     & ~rob_info_3_op1_ready & rob_info_3_is_init & _T_21 ? io_wb_info_i_3_bits_data : _GEN_1604; // @[Rob.scala 269:177 Rob.scala 270:30]
  wire [31:0] _GEN_1610 = io_wb_info_i_3_valid & io_wb_info_i_3_bits_rob_idx == rob_info_3_op2_tag & rob_info_3_is_valid
     & ~rob_info_3_op2_ready & rob_info_3_is_init & _T_21 ? io_wb_info_i_3_bits_data : _GEN_1606; // @[Rob.scala 273:177 Rob.scala 274:30]
  wire [31:0] _GEN_1612 = io_wb_info_i_4_valid & io_wb_info_i_4_bits_rob_idx == rob_info_3_op1_tag & rob_info_3_is_valid
     & ~rob_info_3_op1_ready & rob_info_3_is_init & _T_21 ? io_wb_info_i_4_bits_data : _GEN_1608; // @[Rob.scala 269:177 Rob.scala 270:30]
  wire  _GEN_1613 = io_wb_info_i_4_valid & io_wb_info_i_4_bits_rob_idx == rob_info_3_op1_tag & rob_info_3_is_valid & ~
    rob_info_3_op1_ready & rob_info_3_is_init & _T_21 | (io_wb_info_i_3_valid & io_wb_info_i_3_bits_rob_idx ==
    rob_info_3_op1_tag & rob_info_3_is_valid & ~rob_info_3_op1_ready & rob_info_3_is_init & _T_21 | _GEN_1605); // @[Rob.scala 269:177 Rob.scala 271:31]
  wire [31:0] _GEN_1614 = io_wb_info_i_4_valid & io_wb_info_i_4_bits_rob_idx == rob_info_3_op2_tag & rob_info_3_is_valid
     & ~rob_info_3_op2_ready & rob_info_3_is_init & _T_21 ? io_wb_info_i_4_bits_data : _GEN_1610; // @[Rob.scala 273:177 Rob.scala 274:30]
  wire  _GEN_1615 = io_wb_info_i_4_valid & io_wb_info_i_4_bits_rob_idx == rob_info_3_op2_tag & rob_info_3_is_valid & ~
    rob_info_3_op2_ready & rob_info_3_is_init & _T_21 | (io_wb_info_i_3_valid & io_wb_info_i_3_bits_rob_idx ==
    rob_info_3_op2_tag & rob_info_3_is_valid & ~rob_info_3_op2_ready & rob_info_3_is_init & _T_21 | _GEN_1607); // @[Rob.scala 273:177 Rob.scala 275:31]
  wire [31:0] _GEN_1616 = io_wb_info_i_0_valid & io_wb_info_i_0_bits_rob_idx == rob_info_4_op1_tag & rob_info_4_is_valid
     & ~rob_info_4_op1_ready & rob_info_4_is_init & _T_21 ? io_wb_info_i_0_bits_data : rob_info_4_op1_data; // @[Rob.scala 269:177 Rob.scala 270:30 Rob.scala 175:27]
  wire [31:0] _GEN_1618 = io_wb_info_i_0_valid & io_wb_info_i_0_bits_rob_idx == rob_info_4_op2_tag & rob_info_4_is_valid
     & ~rob_info_4_op2_ready & rob_info_4_is_init & _T_21 ? io_wb_info_i_0_bits_data : rob_info_4_op2_data; // @[Rob.scala 273:177 Rob.scala 274:30 Rob.scala 175:27]
  wire [31:0] _GEN_1620 = io_wb_info_i_1_valid & io_wb_info_i_1_bits_rob_idx == rob_info_4_op1_tag & rob_info_4_is_valid
     & ~rob_info_4_op1_ready & rob_info_4_is_init & _T_21 ? io_wb_info_i_1_bits_data : _GEN_1616; // @[Rob.scala 269:177 Rob.scala 270:30]
  wire [31:0] _GEN_1622 = io_wb_info_i_1_valid & io_wb_info_i_1_bits_rob_idx == rob_info_4_op2_tag & rob_info_4_is_valid
     & ~rob_info_4_op2_ready & rob_info_4_is_init & _T_21 ? io_wb_info_i_1_bits_data : _GEN_1618; // @[Rob.scala 273:177 Rob.scala 274:30]
  wire [31:0] _GEN_1624 = io_wb_info_i_2_valid & io_wb_info_i_2_bits_rob_idx == rob_info_4_op1_tag & rob_info_4_is_valid
     & ~rob_info_4_op1_ready & rob_info_4_is_init & _T_21 ? io_wb_info_i_2_bits_data : _GEN_1620; // @[Rob.scala 269:177 Rob.scala 270:30]
  wire  _GEN_1625 = io_wb_info_i_2_valid & io_wb_info_i_2_bits_rob_idx == rob_info_4_op1_tag & rob_info_4_is_valid & ~
    rob_info_4_op1_ready & rob_info_4_is_init & _T_21 | (io_wb_info_i_1_valid & io_wb_info_i_1_bits_rob_idx ==
    rob_info_4_op1_tag & rob_info_4_is_valid & ~rob_info_4_op1_ready & rob_info_4_is_init & _T_21 | (
    io_wb_info_i_0_valid & io_wb_info_i_0_bits_rob_idx == rob_info_4_op1_tag & rob_info_4_is_valid & ~
    rob_info_4_op1_ready & rob_info_4_is_init & _T_21 | _GEN_1396)); // @[Rob.scala 269:177 Rob.scala 271:31]
  wire [31:0] _GEN_1626 = io_wb_info_i_2_valid & io_wb_info_i_2_bits_rob_idx == rob_info_4_op2_tag & rob_info_4_is_valid
     & ~rob_info_4_op2_ready & rob_info_4_is_init & _T_21 ? io_wb_info_i_2_bits_data : _GEN_1622; // @[Rob.scala 273:177 Rob.scala 274:30]
  wire  _GEN_1627 = io_wb_info_i_2_valid & io_wb_info_i_2_bits_rob_idx == rob_info_4_op2_tag & rob_info_4_is_valid & ~
    rob_info_4_op2_ready & rob_info_4_is_init & _T_21 | (io_wb_info_i_1_valid & io_wb_info_i_1_bits_rob_idx ==
    rob_info_4_op2_tag & rob_info_4_is_valid & ~rob_info_4_op2_ready & rob_info_4_is_init & _T_21 | (
    io_wb_info_i_0_valid & io_wb_info_i_0_bits_rob_idx == rob_info_4_op2_tag & rob_info_4_is_valid & ~
    rob_info_4_op2_ready & rob_info_4_is_init & _T_21 | _GEN_1404)); // @[Rob.scala 273:177 Rob.scala 275:31]
  wire [31:0] _GEN_1628 = io_wb_info_i_3_valid & io_wb_info_i_3_bits_rob_idx == rob_info_4_op1_tag & rob_info_4_is_valid
     & ~rob_info_4_op1_ready & rob_info_4_is_init & _T_21 ? io_wb_info_i_3_bits_data : _GEN_1624; // @[Rob.scala 269:177 Rob.scala 270:30]
  wire [31:0] _GEN_1630 = io_wb_info_i_3_valid & io_wb_info_i_3_bits_rob_idx == rob_info_4_op2_tag & rob_info_4_is_valid
     & ~rob_info_4_op2_ready & rob_info_4_is_init & _T_21 ? io_wb_info_i_3_bits_data : _GEN_1626; // @[Rob.scala 273:177 Rob.scala 274:30]
  wire [31:0] _GEN_1632 = io_wb_info_i_4_valid & io_wb_info_i_4_bits_rob_idx == rob_info_4_op1_tag & rob_info_4_is_valid
     & ~rob_info_4_op1_ready & rob_info_4_is_init & _T_21 ? io_wb_info_i_4_bits_data : _GEN_1628; // @[Rob.scala 269:177 Rob.scala 270:30]
  wire  _GEN_1633 = io_wb_info_i_4_valid & io_wb_info_i_4_bits_rob_idx == rob_info_4_op1_tag & rob_info_4_is_valid & ~
    rob_info_4_op1_ready & rob_info_4_is_init & _T_21 | (io_wb_info_i_3_valid & io_wb_info_i_3_bits_rob_idx ==
    rob_info_4_op1_tag & rob_info_4_is_valid & ~rob_info_4_op1_ready & rob_info_4_is_init & _T_21 | _GEN_1625); // @[Rob.scala 269:177 Rob.scala 271:31]
  wire [31:0] _GEN_1634 = io_wb_info_i_4_valid & io_wb_info_i_4_bits_rob_idx == rob_info_4_op2_tag & rob_info_4_is_valid
     & ~rob_info_4_op2_ready & rob_info_4_is_init & _T_21 ? io_wb_info_i_4_bits_data : _GEN_1630; // @[Rob.scala 273:177 Rob.scala 274:30]
  wire  _GEN_1635 = io_wb_info_i_4_valid & io_wb_info_i_4_bits_rob_idx == rob_info_4_op2_tag & rob_info_4_is_valid & ~
    rob_info_4_op2_ready & rob_info_4_is_init & _T_21 | (io_wb_info_i_3_valid & io_wb_info_i_3_bits_rob_idx ==
    rob_info_4_op2_tag & rob_info_4_is_valid & ~rob_info_4_op2_ready & rob_info_4_is_init & _T_21 | _GEN_1627); // @[Rob.scala 273:177 Rob.scala 275:31]
  wire [31:0] _GEN_1636 = io_wb_info_i_0_valid & io_wb_info_i_0_bits_rob_idx == rob_info_5_op1_tag & rob_info_5_is_valid
     & ~rob_info_5_op1_ready & rob_info_5_is_init & _T_21 ? io_wb_info_i_0_bits_data : rob_info_5_op1_data; // @[Rob.scala 269:177 Rob.scala 270:30 Rob.scala 175:27]
  wire [31:0] _GEN_1638 = io_wb_info_i_0_valid & io_wb_info_i_0_bits_rob_idx == rob_info_5_op2_tag & rob_info_5_is_valid
     & ~rob_info_5_op2_ready & rob_info_5_is_init & _T_21 ? io_wb_info_i_0_bits_data : rob_info_5_op2_data; // @[Rob.scala 273:177 Rob.scala 274:30 Rob.scala 175:27]
  wire [31:0] _GEN_1640 = io_wb_info_i_1_valid & io_wb_info_i_1_bits_rob_idx == rob_info_5_op1_tag & rob_info_5_is_valid
     & ~rob_info_5_op1_ready & rob_info_5_is_init & _T_21 ? io_wb_info_i_1_bits_data : _GEN_1636; // @[Rob.scala 269:177 Rob.scala 270:30]
  wire [31:0] _GEN_1642 = io_wb_info_i_1_valid & io_wb_info_i_1_bits_rob_idx == rob_info_5_op2_tag & rob_info_5_is_valid
     & ~rob_info_5_op2_ready & rob_info_5_is_init & _T_21 ? io_wb_info_i_1_bits_data : _GEN_1638; // @[Rob.scala 273:177 Rob.scala 274:30]
  wire [31:0] _GEN_1644 = io_wb_info_i_2_valid & io_wb_info_i_2_bits_rob_idx == rob_info_5_op1_tag & rob_info_5_is_valid
     & ~rob_info_5_op1_ready & rob_info_5_is_init & _T_21 ? io_wb_info_i_2_bits_data : _GEN_1640; // @[Rob.scala 269:177 Rob.scala 270:30]
  wire  _GEN_1645 = io_wb_info_i_2_valid & io_wb_info_i_2_bits_rob_idx == rob_info_5_op1_tag & rob_info_5_is_valid & ~
    rob_info_5_op1_ready & rob_info_5_is_init & _T_21 | (io_wb_info_i_1_valid & io_wb_info_i_1_bits_rob_idx ==
    rob_info_5_op1_tag & rob_info_5_is_valid & ~rob_info_5_op1_ready & rob_info_5_is_init & _T_21 | (
    io_wb_info_i_0_valid & io_wb_info_i_0_bits_rob_idx == rob_info_5_op1_tag & rob_info_5_is_valid & ~
    rob_info_5_op1_ready & rob_info_5_is_init & _T_21 | _GEN_1397)); // @[Rob.scala 269:177 Rob.scala 271:31]
  wire [31:0] _GEN_1646 = io_wb_info_i_2_valid & io_wb_info_i_2_bits_rob_idx == rob_info_5_op2_tag & rob_info_5_is_valid
     & ~rob_info_5_op2_ready & rob_info_5_is_init & _T_21 ? io_wb_info_i_2_bits_data : _GEN_1642; // @[Rob.scala 273:177 Rob.scala 274:30]
  wire  _GEN_1647 = io_wb_info_i_2_valid & io_wb_info_i_2_bits_rob_idx == rob_info_5_op2_tag & rob_info_5_is_valid & ~
    rob_info_5_op2_ready & rob_info_5_is_init & _T_21 | (io_wb_info_i_1_valid & io_wb_info_i_1_bits_rob_idx ==
    rob_info_5_op2_tag & rob_info_5_is_valid & ~rob_info_5_op2_ready & rob_info_5_is_init & _T_21 | (
    io_wb_info_i_0_valid & io_wb_info_i_0_bits_rob_idx == rob_info_5_op2_tag & rob_info_5_is_valid & ~
    rob_info_5_op2_ready & rob_info_5_is_init & _T_21 | _GEN_1405)); // @[Rob.scala 273:177 Rob.scala 275:31]
  wire [31:0] _GEN_1648 = io_wb_info_i_3_valid & io_wb_info_i_3_bits_rob_idx == rob_info_5_op1_tag & rob_info_5_is_valid
     & ~rob_info_5_op1_ready & rob_info_5_is_init & _T_21 ? io_wb_info_i_3_bits_data : _GEN_1644; // @[Rob.scala 269:177 Rob.scala 270:30]
  wire [31:0] _GEN_1650 = io_wb_info_i_3_valid & io_wb_info_i_3_bits_rob_idx == rob_info_5_op2_tag & rob_info_5_is_valid
     & ~rob_info_5_op2_ready & rob_info_5_is_init & _T_21 ? io_wb_info_i_3_bits_data : _GEN_1646; // @[Rob.scala 273:177 Rob.scala 274:30]
  wire [31:0] _GEN_1652 = io_wb_info_i_4_valid & io_wb_info_i_4_bits_rob_idx == rob_info_5_op1_tag & rob_info_5_is_valid
     & ~rob_info_5_op1_ready & rob_info_5_is_init & _T_21 ? io_wb_info_i_4_bits_data : _GEN_1648; // @[Rob.scala 269:177 Rob.scala 270:30]
  wire  _GEN_1653 = io_wb_info_i_4_valid & io_wb_info_i_4_bits_rob_idx == rob_info_5_op1_tag & rob_info_5_is_valid & ~
    rob_info_5_op1_ready & rob_info_5_is_init & _T_21 | (io_wb_info_i_3_valid & io_wb_info_i_3_bits_rob_idx ==
    rob_info_5_op1_tag & rob_info_5_is_valid & ~rob_info_5_op1_ready & rob_info_5_is_init & _T_21 | _GEN_1645); // @[Rob.scala 269:177 Rob.scala 271:31]
  wire [31:0] _GEN_1654 = io_wb_info_i_4_valid & io_wb_info_i_4_bits_rob_idx == rob_info_5_op2_tag & rob_info_5_is_valid
     & ~rob_info_5_op2_ready & rob_info_5_is_init & _T_21 ? io_wb_info_i_4_bits_data : _GEN_1650; // @[Rob.scala 273:177 Rob.scala 274:30]
  wire  _GEN_1655 = io_wb_info_i_4_valid & io_wb_info_i_4_bits_rob_idx == rob_info_5_op2_tag & rob_info_5_is_valid & ~
    rob_info_5_op2_ready & rob_info_5_is_init & _T_21 | (io_wb_info_i_3_valid & io_wb_info_i_3_bits_rob_idx ==
    rob_info_5_op2_tag & rob_info_5_is_valid & ~rob_info_5_op2_ready & rob_info_5_is_init & _T_21 | _GEN_1647); // @[Rob.scala 273:177 Rob.scala 275:31]
  wire [31:0] _GEN_1656 = io_wb_info_i_0_valid & io_wb_info_i_0_bits_rob_idx == rob_info_6_op1_tag & rob_info_6_is_valid
     & ~rob_info_6_op1_ready & rob_info_6_is_init & _T_21 ? io_wb_info_i_0_bits_data : rob_info_6_op1_data; // @[Rob.scala 269:177 Rob.scala 270:30 Rob.scala 175:27]
  wire [31:0] _GEN_1658 = io_wb_info_i_0_valid & io_wb_info_i_0_bits_rob_idx == rob_info_6_op2_tag & rob_info_6_is_valid
     & ~rob_info_6_op2_ready & rob_info_6_is_init & _T_21 ? io_wb_info_i_0_bits_data : rob_info_6_op2_data; // @[Rob.scala 273:177 Rob.scala 274:30 Rob.scala 175:27]
  wire [31:0] _GEN_1660 = io_wb_info_i_1_valid & io_wb_info_i_1_bits_rob_idx == rob_info_6_op1_tag & rob_info_6_is_valid
     & ~rob_info_6_op1_ready & rob_info_6_is_init & _T_21 ? io_wb_info_i_1_bits_data : _GEN_1656; // @[Rob.scala 269:177 Rob.scala 270:30]
  wire [31:0] _GEN_1662 = io_wb_info_i_1_valid & io_wb_info_i_1_bits_rob_idx == rob_info_6_op2_tag & rob_info_6_is_valid
     & ~rob_info_6_op2_ready & rob_info_6_is_init & _T_21 ? io_wb_info_i_1_bits_data : _GEN_1658; // @[Rob.scala 273:177 Rob.scala 274:30]
  wire [31:0] _GEN_1664 = io_wb_info_i_2_valid & io_wb_info_i_2_bits_rob_idx == rob_info_6_op1_tag & rob_info_6_is_valid
     & ~rob_info_6_op1_ready & rob_info_6_is_init & _T_21 ? io_wb_info_i_2_bits_data : _GEN_1660; // @[Rob.scala 269:177 Rob.scala 270:30]
  wire  _GEN_1665 = io_wb_info_i_2_valid & io_wb_info_i_2_bits_rob_idx == rob_info_6_op1_tag & rob_info_6_is_valid & ~
    rob_info_6_op1_ready & rob_info_6_is_init & _T_21 | (io_wb_info_i_1_valid & io_wb_info_i_1_bits_rob_idx ==
    rob_info_6_op1_tag & rob_info_6_is_valid & ~rob_info_6_op1_ready & rob_info_6_is_init & _T_21 | (
    io_wb_info_i_0_valid & io_wb_info_i_0_bits_rob_idx == rob_info_6_op1_tag & rob_info_6_is_valid & ~
    rob_info_6_op1_ready & rob_info_6_is_init & _T_21 | _GEN_1398)); // @[Rob.scala 269:177 Rob.scala 271:31]
  wire [31:0] _GEN_1666 = io_wb_info_i_2_valid & io_wb_info_i_2_bits_rob_idx == rob_info_6_op2_tag & rob_info_6_is_valid
     & ~rob_info_6_op2_ready & rob_info_6_is_init & _T_21 ? io_wb_info_i_2_bits_data : _GEN_1662; // @[Rob.scala 273:177 Rob.scala 274:30]
  wire  _GEN_1667 = io_wb_info_i_2_valid & io_wb_info_i_2_bits_rob_idx == rob_info_6_op2_tag & rob_info_6_is_valid & ~
    rob_info_6_op2_ready & rob_info_6_is_init & _T_21 | (io_wb_info_i_1_valid & io_wb_info_i_1_bits_rob_idx ==
    rob_info_6_op2_tag & rob_info_6_is_valid & ~rob_info_6_op2_ready & rob_info_6_is_init & _T_21 | (
    io_wb_info_i_0_valid & io_wb_info_i_0_bits_rob_idx == rob_info_6_op2_tag & rob_info_6_is_valid & ~
    rob_info_6_op2_ready & rob_info_6_is_init & _T_21 | _GEN_1406)); // @[Rob.scala 273:177 Rob.scala 275:31]
  wire [31:0] _GEN_1668 = io_wb_info_i_3_valid & io_wb_info_i_3_bits_rob_idx == rob_info_6_op1_tag & rob_info_6_is_valid
     & ~rob_info_6_op1_ready & rob_info_6_is_init & _T_21 ? io_wb_info_i_3_bits_data : _GEN_1664; // @[Rob.scala 269:177 Rob.scala 270:30]
  wire [31:0] _GEN_1670 = io_wb_info_i_3_valid & io_wb_info_i_3_bits_rob_idx == rob_info_6_op2_tag & rob_info_6_is_valid
     & ~rob_info_6_op2_ready & rob_info_6_is_init & _T_21 ? io_wb_info_i_3_bits_data : _GEN_1666; // @[Rob.scala 273:177 Rob.scala 274:30]
  wire [31:0] _GEN_1672 = io_wb_info_i_4_valid & io_wb_info_i_4_bits_rob_idx == rob_info_6_op1_tag & rob_info_6_is_valid
     & ~rob_info_6_op1_ready & rob_info_6_is_init & _T_21 ? io_wb_info_i_4_bits_data : _GEN_1668; // @[Rob.scala 269:177 Rob.scala 270:30]
  wire  _GEN_1673 = io_wb_info_i_4_valid & io_wb_info_i_4_bits_rob_idx == rob_info_6_op1_tag & rob_info_6_is_valid & ~
    rob_info_6_op1_ready & rob_info_6_is_init & _T_21 | (io_wb_info_i_3_valid & io_wb_info_i_3_bits_rob_idx ==
    rob_info_6_op1_tag & rob_info_6_is_valid & ~rob_info_6_op1_ready & rob_info_6_is_init & _T_21 | _GEN_1665); // @[Rob.scala 269:177 Rob.scala 271:31]
  wire [31:0] _GEN_1674 = io_wb_info_i_4_valid & io_wb_info_i_4_bits_rob_idx == rob_info_6_op2_tag & rob_info_6_is_valid
     & ~rob_info_6_op2_ready & rob_info_6_is_init & _T_21 ? io_wb_info_i_4_bits_data : _GEN_1670; // @[Rob.scala 273:177 Rob.scala 274:30]
  wire  _GEN_1675 = io_wb_info_i_4_valid & io_wb_info_i_4_bits_rob_idx == rob_info_6_op2_tag & rob_info_6_is_valid & ~
    rob_info_6_op2_ready & rob_info_6_is_init & _T_21 | (io_wb_info_i_3_valid & io_wb_info_i_3_bits_rob_idx ==
    rob_info_6_op2_tag & rob_info_6_is_valid & ~rob_info_6_op2_ready & rob_info_6_is_init & _T_21 | _GEN_1667); // @[Rob.scala 273:177 Rob.scala 275:31]
  wire [31:0] _GEN_1676 = io_wb_info_i_0_valid & io_wb_info_i_0_bits_rob_idx == rob_info_7_op1_tag & rob_info_7_is_valid
     & ~rob_info_7_op1_ready & rob_info_7_is_init & _T_21 ? io_wb_info_i_0_bits_data : rob_info_7_op1_data; // @[Rob.scala 269:177 Rob.scala 270:30 Rob.scala 175:27]
  wire [31:0] _GEN_1678 = io_wb_info_i_0_valid & io_wb_info_i_0_bits_rob_idx == rob_info_7_op2_tag & rob_info_7_is_valid
     & ~rob_info_7_op2_ready & rob_info_7_is_init & _T_21 ? io_wb_info_i_0_bits_data : rob_info_7_op2_data; // @[Rob.scala 273:177 Rob.scala 274:30 Rob.scala 175:27]
  wire [31:0] _GEN_1680 = io_wb_info_i_1_valid & io_wb_info_i_1_bits_rob_idx == rob_info_7_op1_tag & rob_info_7_is_valid
     & ~rob_info_7_op1_ready & rob_info_7_is_init & _T_21 ? io_wb_info_i_1_bits_data : _GEN_1676; // @[Rob.scala 269:177 Rob.scala 270:30]
  wire [31:0] _GEN_1682 = io_wb_info_i_1_valid & io_wb_info_i_1_bits_rob_idx == rob_info_7_op2_tag & rob_info_7_is_valid
     & ~rob_info_7_op2_ready & rob_info_7_is_init & _T_21 ? io_wb_info_i_1_bits_data : _GEN_1678; // @[Rob.scala 273:177 Rob.scala 274:30]
  wire [31:0] _GEN_1684 = io_wb_info_i_2_valid & io_wb_info_i_2_bits_rob_idx == rob_info_7_op1_tag & rob_info_7_is_valid
     & ~rob_info_7_op1_ready & rob_info_7_is_init & _T_21 ? io_wb_info_i_2_bits_data : _GEN_1680; // @[Rob.scala 269:177 Rob.scala 270:30]
  wire  _GEN_1685 = io_wb_info_i_2_valid & io_wb_info_i_2_bits_rob_idx == rob_info_7_op1_tag & rob_info_7_is_valid & ~
    rob_info_7_op1_ready & rob_info_7_is_init & _T_21 | (io_wb_info_i_1_valid & io_wb_info_i_1_bits_rob_idx ==
    rob_info_7_op1_tag & rob_info_7_is_valid & ~rob_info_7_op1_ready & rob_info_7_is_init & _T_21 | (
    io_wb_info_i_0_valid & io_wb_info_i_0_bits_rob_idx == rob_info_7_op1_tag & rob_info_7_is_valid & ~
    rob_info_7_op1_ready & rob_info_7_is_init & _T_21 | _GEN_1399)); // @[Rob.scala 269:177 Rob.scala 271:31]
  wire [31:0] _GEN_1686 = io_wb_info_i_2_valid & io_wb_info_i_2_bits_rob_idx == rob_info_7_op2_tag & rob_info_7_is_valid
     & ~rob_info_7_op2_ready & rob_info_7_is_init & _T_21 ? io_wb_info_i_2_bits_data : _GEN_1682; // @[Rob.scala 273:177 Rob.scala 274:30]
  wire  _GEN_1687 = io_wb_info_i_2_valid & io_wb_info_i_2_bits_rob_idx == rob_info_7_op2_tag & rob_info_7_is_valid & ~
    rob_info_7_op2_ready & rob_info_7_is_init & _T_21 | (io_wb_info_i_1_valid & io_wb_info_i_1_bits_rob_idx ==
    rob_info_7_op2_tag & rob_info_7_is_valid & ~rob_info_7_op2_ready & rob_info_7_is_init & _T_21 | (
    io_wb_info_i_0_valid & io_wb_info_i_0_bits_rob_idx == rob_info_7_op2_tag & rob_info_7_is_valid & ~
    rob_info_7_op2_ready & rob_info_7_is_init & _T_21 | _GEN_1407)); // @[Rob.scala 273:177 Rob.scala 275:31]
  wire [31:0] _GEN_1688 = io_wb_info_i_3_valid & io_wb_info_i_3_bits_rob_idx == rob_info_7_op1_tag & rob_info_7_is_valid
     & ~rob_info_7_op1_ready & rob_info_7_is_init & _T_21 ? io_wb_info_i_3_bits_data : _GEN_1684; // @[Rob.scala 269:177 Rob.scala 270:30]
  wire [31:0] _GEN_1690 = io_wb_info_i_3_valid & io_wb_info_i_3_bits_rob_idx == rob_info_7_op2_tag & rob_info_7_is_valid
     & ~rob_info_7_op2_ready & rob_info_7_is_init & _T_21 ? io_wb_info_i_3_bits_data : _GEN_1686; // @[Rob.scala 273:177 Rob.scala 274:30]
  wire [31:0] _GEN_1692 = io_wb_info_i_4_valid & io_wb_info_i_4_bits_rob_idx == rob_info_7_op1_tag & rob_info_7_is_valid
     & ~rob_info_7_op1_ready & rob_info_7_is_init & _T_21 ? io_wb_info_i_4_bits_data : _GEN_1688; // @[Rob.scala 269:177 Rob.scala 270:30]
  wire  _GEN_1693 = io_wb_info_i_4_valid & io_wb_info_i_4_bits_rob_idx == rob_info_7_op1_tag & rob_info_7_is_valid & ~
    rob_info_7_op1_ready & rob_info_7_is_init & _T_21 | (io_wb_info_i_3_valid & io_wb_info_i_3_bits_rob_idx ==
    rob_info_7_op1_tag & rob_info_7_is_valid & ~rob_info_7_op1_ready & rob_info_7_is_init & _T_21 | _GEN_1685); // @[Rob.scala 269:177 Rob.scala 271:31]
  wire [31:0] _GEN_1694 = io_wb_info_i_4_valid & io_wb_info_i_4_bits_rob_idx == rob_info_7_op2_tag & rob_info_7_is_valid
     & ~rob_info_7_op2_ready & rob_info_7_is_init & _T_21 ? io_wb_info_i_4_bits_data : _GEN_1690; // @[Rob.scala 273:177 Rob.scala 274:30]
  wire  _GEN_1695 = io_wb_info_i_4_valid & io_wb_info_i_4_bits_rob_idx == rob_info_7_op2_tag & rob_info_7_is_valid & ~
    rob_info_7_op2_ready & rob_info_7_is_init & _T_21 | (io_wb_info_i_3_valid & io_wb_info_i_3_bits_rob_idx ==
    rob_info_7_op2_tag & rob_info_7_is_valid & ~rob_info_7_op2_ready & rob_info_7_is_init & _T_21 | _GEN_1687); // @[Rob.scala 273:177 Rob.scala 275:31]
  wire  _GEN_1697 = 3'h1 == io_wb_info_i_0_bits_rob_idx ? rob_info_1_is_valid : rob_info_0_is_valid; // @[Rob.scala 283:31 Rob.scala 283:31]
  wire  _GEN_1698 = 3'h2 == io_wb_info_i_0_bits_rob_idx ? rob_info_2_is_valid : _GEN_1697; // @[Rob.scala 283:31 Rob.scala 283:31]
  wire  _GEN_1699 = 3'h3 == io_wb_info_i_0_bits_rob_idx ? rob_info_3_is_valid : _GEN_1698; // @[Rob.scala 283:31 Rob.scala 283:31]
  wire  _GEN_1700 = 3'h4 == io_wb_info_i_0_bits_rob_idx ? rob_info_4_is_valid : _GEN_1699; // @[Rob.scala 283:31 Rob.scala 283:31]
  wire  _GEN_1701 = 3'h5 == io_wb_info_i_0_bits_rob_idx ? rob_info_5_is_valid : _GEN_1700; // @[Rob.scala 283:31 Rob.scala 283:31]
  wire  _GEN_1702 = 3'h6 == io_wb_info_i_0_bits_rob_idx ? rob_info_6_is_valid : _GEN_1701; // @[Rob.scala 283:31 Rob.scala 283:31]
  wire  _GEN_1703 = 3'h7 == io_wb_info_i_0_bits_rob_idx ? rob_info_7_is_valid : _GEN_1702; // @[Rob.scala 283:31 Rob.scala 283:31]
  wire [31:0] _GEN_1704 = 3'h0 == io_wb_info_i_0_bits_rob_idx ? io_wb_info_i_0_bits_data : rob_info_0_commit_data; // @[Rob.scala 284:37 Rob.scala 284:37 Rob.scala 175:27]
  wire [31:0] _GEN_1705 = 3'h1 == io_wb_info_i_0_bits_rob_idx ? io_wb_info_i_0_bits_data : rob_info_1_commit_data; // @[Rob.scala 284:37 Rob.scala 284:37 Rob.scala 175:27]
  wire [31:0] _GEN_1706 = 3'h2 == io_wb_info_i_0_bits_rob_idx ? io_wb_info_i_0_bits_data : rob_info_2_commit_data; // @[Rob.scala 284:37 Rob.scala 284:37 Rob.scala 175:27]
  wire [31:0] _GEN_1707 = 3'h3 == io_wb_info_i_0_bits_rob_idx ? io_wb_info_i_0_bits_data : rob_info_3_commit_data; // @[Rob.scala 284:37 Rob.scala 284:37 Rob.scala 175:27]
  wire [31:0] _GEN_1708 = 3'h4 == io_wb_info_i_0_bits_rob_idx ? io_wb_info_i_0_bits_data : rob_info_4_commit_data; // @[Rob.scala 284:37 Rob.scala 284:37 Rob.scala 175:27]
  wire [31:0] _GEN_1709 = 3'h5 == io_wb_info_i_0_bits_rob_idx ? io_wb_info_i_0_bits_data : rob_info_5_commit_data; // @[Rob.scala 284:37 Rob.scala 284:37 Rob.scala 175:27]
  wire [31:0] _GEN_1710 = 3'h6 == io_wb_info_i_0_bits_rob_idx ? io_wb_info_i_0_bits_data : rob_info_6_commit_data; // @[Rob.scala 284:37 Rob.scala 284:37 Rob.scala 175:27]
  wire [31:0] _GEN_1711 = 3'h7 == io_wb_info_i_0_bits_rob_idx ? io_wb_info_i_0_bits_data : rob_info_7_commit_data; // @[Rob.scala 284:37 Rob.scala 284:37 Rob.scala 175:27]
  wire  _GEN_1712 = 3'h0 == io_wb_info_i_0_bits_rob_idx | _GEN_1368; // @[Rob.scala 285:38 Rob.scala 285:38]
  wire  _GEN_1713 = 3'h1 == io_wb_info_i_0_bits_rob_idx | _GEN_1369; // @[Rob.scala 285:38 Rob.scala 285:38]
  wire  _GEN_1714 = 3'h2 == io_wb_info_i_0_bits_rob_idx | _GEN_1370; // @[Rob.scala 285:38 Rob.scala 285:38]
  wire  _GEN_1715 = 3'h3 == io_wb_info_i_0_bits_rob_idx | _GEN_1371; // @[Rob.scala 285:38 Rob.scala 285:38]
  wire  _GEN_1716 = 3'h4 == io_wb_info_i_0_bits_rob_idx | _GEN_1372; // @[Rob.scala 285:38 Rob.scala 285:38]
  wire  _GEN_1717 = 3'h5 == io_wb_info_i_0_bits_rob_idx | _GEN_1373; // @[Rob.scala 285:38 Rob.scala 285:38]
  wire  _GEN_1718 = 3'h6 == io_wb_info_i_0_bits_rob_idx | _GEN_1374; // @[Rob.scala 285:38 Rob.scala 285:38]
  wire  _GEN_1719 = 3'h7 == io_wb_info_i_0_bits_rob_idx | _GEN_1375; // @[Rob.scala 285:38 Rob.scala 285:38]
  wire  _GEN_1720 = 3'h0 == io_wb_info_i_0_bits_rob_idx ? 1'h0 : _GEN_1376; // @[Rob.scala 286:30 Rob.scala 286:30]
  wire  _GEN_1721 = 3'h1 == io_wb_info_i_0_bits_rob_idx ? 1'h0 : _GEN_1377; // @[Rob.scala 286:30 Rob.scala 286:30]
  wire  _GEN_1722 = 3'h2 == io_wb_info_i_0_bits_rob_idx ? 1'h0 : _GEN_1378; // @[Rob.scala 286:30 Rob.scala 286:30]
  wire  _GEN_1723 = 3'h3 == io_wb_info_i_0_bits_rob_idx ? 1'h0 : _GEN_1379; // @[Rob.scala 286:30 Rob.scala 286:30]
  wire  _GEN_1724 = 3'h4 == io_wb_info_i_0_bits_rob_idx ? 1'h0 : _GEN_1380; // @[Rob.scala 286:30 Rob.scala 286:30]
  wire  _GEN_1725 = 3'h5 == io_wb_info_i_0_bits_rob_idx ? 1'h0 : _GEN_1381; // @[Rob.scala 286:30 Rob.scala 286:30]
  wire  _GEN_1726 = 3'h6 == io_wb_info_i_0_bits_rob_idx ? 1'h0 : _GEN_1382; // @[Rob.scala 286:30 Rob.scala 286:30]
  wire  _GEN_1727 = 3'h7 == io_wb_info_i_0_bits_rob_idx ? 1'h0 : _GEN_1383; // @[Rob.scala 286:30 Rob.scala 286:30]
  wire  _GEN_1728 = 3'h0 == io_wb_info_i_0_bits_rob_idx ? 1'h0 : _GEN_1416; // @[Rob.scala 287:34 Rob.scala 287:34]
  wire  _GEN_1729 = 3'h1 == io_wb_info_i_0_bits_rob_idx ? 1'h0 : _GEN_1417; // @[Rob.scala 287:34 Rob.scala 287:34]
  wire  _GEN_1730 = 3'h2 == io_wb_info_i_0_bits_rob_idx ? 1'h0 : _GEN_1418; // @[Rob.scala 287:34 Rob.scala 287:34]
  wire  _GEN_1731 = 3'h3 == io_wb_info_i_0_bits_rob_idx ? 1'h0 : _GEN_1419; // @[Rob.scala 287:34 Rob.scala 287:34]
  wire  _GEN_1732 = 3'h4 == io_wb_info_i_0_bits_rob_idx ? 1'h0 : _GEN_1420; // @[Rob.scala 287:34 Rob.scala 287:34]
  wire  _GEN_1733 = 3'h5 == io_wb_info_i_0_bits_rob_idx ? 1'h0 : _GEN_1421; // @[Rob.scala 287:34 Rob.scala 287:34]
  wire  _GEN_1734 = 3'h6 == io_wb_info_i_0_bits_rob_idx ? 1'h0 : _GEN_1422; // @[Rob.scala 287:34 Rob.scala 287:34]
  wire  _GEN_1735 = 3'h7 == io_wb_info_i_0_bits_rob_idx ? 1'h0 : _GEN_1423; // @[Rob.scala 287:34 Rob.scala 287:34]
  wire  _GEN_1736 = 3'h0 == io_wb_info_i_0_bits_rob_idx ? 1'h0 : _GEN_1408; // @[Rob.scala 288:38 Rob.scala 288:38]
  wire  _GEN_1737 = 3'h1 == io_wb_info_i_0_bits_rob_idx ? 1'h0 : _GEN_1409; // @[Rob.scala 288:38 Rob.scala 288:38]
  wire  _GEN_1738 = 3'h2 == io_wb_info_i_0_bits_rob_idx ? 1'h0 : _GEN_1410; // @[Rob.scala 288:38 Rob.scala 288:38]
  wire  _GEN_1739 = 3'h3 == io_wb_info_i_0_bits_rob_idx ? 1'h0 : _GEN_1411; // @[Rob.scala 288:38 Rob.scala 288:38]
  wire  _GEN_1740 = 3'h4 == io_wb_info_i_0_bits_rob_idx ? 1'h0 : _GEN_1412; // @[Rob.scala 288:38 Rob.scala 288:38]
  wire  _GEN_1741 = 3'h5 == io_wb_info_i_0_bits_rob_idx ? 1'h0 : _GEN_1413; // @[Rob.scala 288:38 Rob.scala 288:38]
  wire  _GEN_1742 = 3'h6 == io_wb_info_i_0_bits_rob_idx ? 1'h0 : _GEN_1414; // @[Rob.scala 288:38 Rob.scala 288:38]
  wire  _GEN_1743 = 3'h7 == io_wb_info_i_0_bits_rob_idx ? 1'h0 : _GEN_1415; // @[Rob.scala 288:38 Rob.scala 288:38]
  wire [31:0] _GEN_1744 = 3'h0 == io_wb_info_i_0_bits_rob_idx ? 32'h0 : _GEN_1512; // @[Rob.scala 289:34 Rob.scala 289:34]
  wire [31:0] _GEN_1745 = 3'h1 == io_wb_info_i_0_bits_rob_idx ? 32'h0 : _GEN_1513; // @[Rob.scala 289:34 Rob.scala 289:34]
  wire [31:0] _GEN_1746 = 3'h2 == io_wb_info_i_0_bits_rob_idx ? 32'h0 : _GEN_1514; // @[Rob.scala 289:34 Rob.scala 289:34]
  wire [31:0] _GEN_1747 = 3'h3 == io_wb_info_i_0_bits_rob_idx ? 32'h0 : _GEN_1515; // @[Rob.scala 289:34 Rob.scala 289:34]
  wire [31:0] _GEN_1748 = 3'h4 == io_wb_info_i_0_bits_rob_idx ? 32'h0 : _GEN_1516; // @[Rob.scala 289:34 Rob.scala 289:34]
  wire [31:0] _GEN_1749 = 3'h5 == io_wb_info_i_0_bits_rob_idx ? 32'h0 : _GEN_1517; // @[Rob.scala 289:34 Rob.scala 289:34]
  wire [31:0] _GEN_1750 = 3'h6 == io_wb_info_i_0_bits_rob_idx ? 32'h0 : _GEN_1518; // @[Rob.scala 289:34 Rob.scala 289:34]
  wire [31:0] _GEN_1751 = 3'h7 == io_wb_info_i_0_bits_rob_idx ? 32'h0 : _GEN_1519; // @[Rob.scala 289:34 Rob.scala 289:34]
  wire [31:0] _GEN_1752 = io_wb_info_i_0_valid & _GEN_1703 & _T_21 ? _GEN_1704 : rob_info_0_commit_data; // @[Rob.scala 283:75 Rob.scala 175:27]
  wire [31:0] _GEN_1753 = io_wb_info_i_0_valid & _GEN_1703 & _T_21 ? _GEN_1705 : rob_info_1_commit_data; // @[Rob.scala 283:75 Rob.scala 175:27]
  wire [31:0] _GEN_1754 = io_wb_info_i_0_valid & _GEN_1703 & _T_21 ? _GEN_1706 : rob_info_2_commit_data; // @[Rob.scala 283:75 Rob.scala 175:27]
  wire [31:0] _GEN_1755 = io_wb_info_i_0_valid & _GEN_1703 & _T_21 ? _GEN_1707 : rob_info_3_commit_data; // @[Rob.scala 283:75 Rob.scala 175:27]
  wire [31:0] _GEN_1756 = io_wb_info_i_0_valid & _GEN_1703 & _T_21 ? _GEN_1708 : rob_info_4_commit_data; // @[Rob.scala 283:75 Rob.scala 175:27]
  wire [31:0] _GEN_1757 = io_wb_info_i_0_valid & _GEN_1703 & _T_21 ? _GEN_1709 : rob_info_5_commit_data; // @[Rob.scala 283:75 Rob.scala 175:27]
  wire [31:0] _GEN_1758 = io_wb_info_i_0_valid & _GEN_1703 & _T_21 ? _GEN_1710 : rob_info_6_commit_data; // @[Rob.scala 283:75 Rob.scala 175:27]
  wire [31:0] _GEN_1759 = io_wb_info_i_0_valid & _GEN_1703 & _T_21 ? _GEN_1711 : rob_info_7_commit_data; // @[Rob.scala 283:75 Rob.scala 175:27]
  wire  _GEN_1760 = io_wb_info_i_0_valid & _GEN_1703 & _T_21 ? _GEN_1712 : _GEN_1368; // @[Rob.scala 283:75]
  wire  _GEN_1761 = io_wb_info_i_0_valid & _GEN_1703 & _T_21 ? _GEN_1713 : _GEN_1369; // @[Rob.scala 283:75]
  wire  _GEN_1762 = io_wb_info_i_0_valid & _GEN_1703 & _T_21 ? _GEN_1714 : _GEN_1370; // @[Rob.scala 283:75]
  wire  _GEN_1763 = io_wb_info_i_0_valid & _GEN_1703 & _T_21 ? _GEN_1715 : _GEN_1371; // @[Rob.scala 283:75]
  wire  _GEN_1764 = io_wb_info_i_0_valid & _GEN_1703 & _T_21 ? _GEN_1716 : _GEN_1372; // @[Rob.scala 283:75]
  wire  _GEN_1765 = io_wb_info_i_0_valid & _GEN_1703 & _T_21 ? _GEN_1717 : _GEN_1373; // @[Rob.scala 283:75]
  wire  _GEN_1766 = io_wb_info_i_0_valid & _GEN_1703 & _T_21 ? _GEN_1718 : _GEN_1374; // @[Rob.scala 283:75]
  wire  _GEN_1767 = io_wb_info_i_0_valid & _GEN_1703 & _T_21 ? _GEN_1719 : _GEN_1375; // @[Rob.scala 283:75]
  wire  _GEN_1768 = io_wb_info_i_0_valid & _GEN_1703 & _T_21 ? _GEN_1720 : _GEN_1376; // @[Rob.scala 283:75]
  wire  _GEN_1769 = io_wb_info_i_0_valid & _GEN_1703 & _T_21 ? _GEN_1721 : _GEN_1377; // @[Rob.scala 283:75]
  wire  _GEN_1770 = io_wb_info_i_0_valid & _GEN_1703 & _T_21 ? _GEN_1722 : _GEN_1378; // @[Rob.scala 283:75]
  wire  _GEN_1771 = io_wb_info_i_0_valid & _GEN_1703 & _T_21 ? _GEN_1723 : _GEN_1379; // @[Rob.scala 283:75]
  wire  _GEN_1772 = io_wb_info_i_0_valid & _GEN_1703 & _T_21 ? _GEN_1724 : _GEN_1380; // @[Rob.scala 283:75]
  wire  _GEN_1773 = io_wb_info_i_0_valid & _GEN_1703 & _T_21 ? _GEN_1725 : _GEN_1381; // @[Rob.scala 283:75]
  wire  _GEN_1774 = io_wb_info_i_0_valid & _GEN_1703 & _T_21 ? _GEN_1726 : _GEN_1382; // @[Rob.scala 283:75]
  wire  _GEN_1775 = io_wb_info_i_0_valid & _GEN_1703 & _T_21 ? _GEN_1727 : _GEN_1383; // @[Rob.scala 283:75]
  wire  _GEN_1776 = io_wb_info_i_0_valid & _GEN_1703 & _T_21 ? _GEN_1728 : _GEN_1416; // @[Rob.scala 283:75]
  wire  _GEN_1777 = io_wb_info_i_0_valid & _GEN_1703 & _T_21 ? _GEN_1729 : _GEN_1417; // @[Rob.scala 283:75]
  wire  _GEN_1778 = io_wb_info_i_0_valid & _GEN_1703 & _T_21 ? _GEN_1730 : _GEN_1418; // @[Rob.scala 283:75]
  wire  _GEN_1779 = io_wb_info_i_0_valid & _GEN_1703 & _T_21 ? _GEN_1731 : _GEN_1419; // @[Rob.scala 283:75]
  wire  _GEN_1780 = io_wb_info_i_0_valid & _GEN_1703 & _T_21 ? _GEN_1732 : _GEN_1420; // @[Rob.scala 283:75]
  wire  _GEN_1781 = io_wb_info_i_0_valid & _GEN_1703 & _T_21 ? _GEN_1733 : _GEN_1421; // @[Rob.scala 283:75]
  wire  _GEN_1782 = io_wb_info_i_0_valid & _GEN_1703 & _T_21 ? _GEN_1734 : _GEN_1422; // @[Rob.scala 283:75]
  wire  _GEN_1783 = io_wb_info_i_0_valid & _GEN_1703 & _T_21 ? _GEN_1735 : _GEN_1423; // @[Rob.scala 283:75]
  wire  _GEN_1784 = io_wb_info_i_0_valid & _GEN_1703 & _T_21 ? _GEN_1736 : _GEN_1408; // @[Rob.scala 283:75]
  wire  _GEN_1785 = io_wb_info_i_0_valid & _GEN_1703 & _T_21 ? _GEN_1737 : _GEN_1409; // @[Rob.scala 283:75]
  wire  _GEN_1786 = io_wb_info_i_0_valid & _GEN_1703 & _T_21 ? _GEN_1738 : _GEN_1410; // @[Rob.scala 283:75]
  wire  _GEN_1787 = io_wb_info_i_0_valid & _GEN_1703 & _T_21 ? _GEN_1739 : _GEN_1411; // @[Rob.scala 283:75]
  wire  _GEN_1788 = io_wb_info_i_0_valid & _GEN_1703 & _T_21 ? _GEN_1740 : _GEN_1412; // @[Rob.scala 283:75]
  wire  _GEN_1789 = io_wb_info_i_0_valid & _GEN_1703 & _T_21 ? _GEN_1741 : _GEN_1413; // @[Rob.scala 283:75]
  wire  _GEN_1790 = io_wb_info_i_0_valid & _GEN_1703 & _T_21 ? _GEN_1742 : _GEN_1414; // @[Rob.scala 283:75]
  wire  _GEN_1791 = io_wb_info_i_0_valid & _GEN_1703 & _T_21 ? _GEN_1743 : _GEN_1415; // @[Rob.scala 283:75]
  wire [31:0] _GEN_1792 = io_wb_info_i_0_valid & _GEN_1703 & _T_21 ? _GEN_1744 : _GEN_1512; // @[Rob.scala 283:75]
  wire [31:0] _GEN_1793 = io_wb_info_i_0_valid & _GEN_1703 & _T_21 ? _GEN_1745 : _GEN_1513; // @[Rob.scala 283:75]
  wire [31:0] _GEN_1794 = io_wb_info_i_0_valid & _GEN_1703 & _T_21 ? _GEN_1746 : _GEN_1514; // @[Rob.scala 283:75]
  wire [31:0] _GEN_1795 = io_wb_info_i_0_valid & _GEN_1703 & _T_21 ? _GEN_1747 : _GEN_1515; // @[Rob.scala 283:75]
  wire [31:0] _GEN_1796 = io_wb_info_i_0_valid & _GEN_1703 & _T_21 ? _GEN_1748 : _GEN_1516; // @[Rob.scala 283:75]
  wire [31:0] _GEN_1797 = io_wb_info_i_0_valid & _GEN_1703 & _T_21 ? _GEN_1749 : _GEN_1517; // @[Rob.scala 283:75]
  wire [31:0] _GEN_1798 = io_wb_info_i_0_valid & _GEN_1703 & _T_21 ? _GEN_1750 : _GEN_1518; // @[Rob.scala 283:75]
  wire [31:0] _GEN_1799 = io_wb_info_i_0_valid & _GEN_1703 & _T_21 ? _GEN_1751 : _GEN_1519; // @[Rob.scala 283:75]
  wire  _GEN_1801 = 3'h1 == io_wb_info_i_1_bits_rob_idx ? rob_info_1_is_valid : rob_info_0_is_valid; // @[Rob.scala 283:31 Rob.scala 283:31]
  wire  _GEN_1802 = 3'h2 == io_wb_info_i_1_bits_rob_idx ? rob_info_2_is_valid : _GEN_1801; // @[Rob.scala 283:31 Rob.scala 283:31]
  wire  _GEN_1803 = 3'h3 == io_wb_info_i_1_bits_rob_idx ? rob_info_3_is_valid : _GEN_1802; // @[Rob.scala 283:31 Rob.scala 283:31]
  wire  _GEN_1804 = 3'h4 == io_wb_info_i_1_bits_rob_idx ? rob_info_4_is_valid : _GEN_1803; // @[Rob.scala 283:31 Rob.scala 283:31]
  wire  _GEN_1805 = 3'h5 == io_wb_info_i_1_bits_rob_idx ? rob_info_5_is_valid : _GEN_1804; // @[Rob.scala 283:31 Rob.scala 283:31]
  wire  _GEN_1806 = 3'h6 == io_wb_info_i_1_bits_rob_idx ? rob_info_6_is_valid : _GEN_1805; // @[Rob.scala 283:31 Rob.scala 283:31]
  wire  _GEN_1807 = 3'h7 == io_wb_info_i_1_bits_rob_idx ? rob_info_7_is_valid : _GEN_1806; // @[Rob.scala 283:31 Rob.scala 283:31]
  wire [31:0] _GEN_1808 = 3'h0 == io_wb_info_i_1_bits_rob_idx ? io_wb_info_i_1_bits_data : _GEN_1752; // @[Rob.scala 284:37 Rob.scala 284:37]
  wire [31:0] _GEN_1809 = 3'h1 == io_wb_info_i_1_bits_rob_idx ? io_wb_info_i_1_bits_data : _GEN_1753; // @[Rob.scala 284:37 Rob.scala 284:37]
  wire [31:0] _GEN_1810 = 3'h2 == io_wb_info_i_1_bits_rob_idx ? io_wb_info_i_1_bits_data : _GEN_1754; // @[Rob.scala 284:37 Rob.scala 284:37]
  wire [31:0] _GEN_1811 = 3'h3 == io_wb_info_i_1_bits_rob_idx ? io_wb_info_i_1_bits_data : _GEN_1755; // @[Rob.scala 284:37 Rob.scala 284:37]
  wire [31:0] _GEN_1812 = 3'h4 == io_wb_info_i_1_bits_rob_idx ? io_wb_info_i_1_bits_data : _GEN_1756; // @[Rob.scala 284:37 Rob.scala 284:37]
  wire [31:0] _GEN_1813 = 3'h5 == io_wb_info_i_1_bits_rob_idx ? io_wb_info_i_1_bits_data : _GEN_1757; // @[Rob.scala 284:37 Rob.scala 284:37]
  wire [31:0] _GEN_1814 = 3'h6 == io_wb_info_i_1_bits_rob_idx ? io_wb_info_i_1_bits_data : _GEN_1758; // @[Rob.scala 284:37 Rob.scala 284:37]
  wire [31:0] _GEN_1815 = 3'h7 == io_wb_info_i_1_bits_rob_idx ? io_wb_info_i_1_bits_data : _GEN_1759; // @[Rob.scala 284:37 Rob.scala 284:37]
  wire  _GEN_1816 = 3'h0 == io_wb_info_i_1_bits_rob_idx | _GEN_1760; // @[Rob.scala 285:38 Rob.scala 285:38]
  wire  _GEN_1817 = 3'h1 == io_wb_info_i_1_bits_rob_idx | _GEN_1761; // @[Rob.scala 285:38 Rob.scala 285:38]
  wire  _GEN_1818 = 3'h2 == io_wb_info_i_1_bits_rob_idx | _GEN_1762; // @[Rob.scala 285:38 Rob.scala 285:38]
  wire  _GEN_1819 = 3'h3 == io_wb_info_i_1_bits_rob_idx | _GEN_1763; // @[Rob.scala 285:38 Rob.scala 285:38]
  wire  _GEN_1820 = 3'h4 == io_wb_info_i_1_bits_rob_idx | _GEN_1764; // @[Rob.scala 285:38 Rob.scala 285:38]
  wire  _GEN_1821 = 3'h5 == io_wb_info_i_1_bits_rob_idx | _GEN_1765; // @[Rob.scala 285:38 Rob.scala 285:38]
  wire  _GEN_1822 = 3'h6 == io_wb_info_i_1_bits_rob_idx | _GEN_1766; // @[Rob.scala 285:38 Rob.scala 285:38]
  wire  _GEN_1823 = 3'h7 == io_wb_info_i_1_bits_rob_idx | _GEN_1767; // @[Rob.scala 285:38 Rob.scala 285:38]
  wire  _GEN_1824 = 3'h0 == io_wb_info_i_1_bits_rob_idx ? 1'h0 : _GEN_1768; // @[Rob.scala 286:30 Rob.scala 286:30]
  wire  _GEN_1825 = 3'h1 == io_wb_info_i_1_bits_rob_idx ? 1'h0 : _GEN_1769; // @[Rob.scala 286:30 Rob.scala 286:30]
  wire  _GEN_1826 = 3'h2 == io_wb_info_i_1_bits_rob_idx ? 1'h0 : _GEN_1770; // @[Rob.scala 286:30 Rob.scala 286:30]
  wire  _GEN_1827 = 3'h3 == io_wb_info_i_1_bits_rob_idx ? 1'h0 : _GEN_1771; // @[Rob.scala 286:30 Rob.scala 286:30]
  wire  _GEN_1828 = 3'h4 == io_wb_info_i_1_bits_rob_idx ? 1'h0 : _GEN_1772; // @[Rob.scala 286:30 Rob.scala 286:30]
  wire  _GEN_1829 = 3'h5 == io_wb_info_i_1_bits_rob_idx ? 1'h0 : _GEN_1773; // @[Rob.scala 286:30 Rob.scala 286:30]
  wire  _GEN_1830 = 3'h6 == io_wb_info_i_1_bits_rob_idx ? 1'h0 : _GEN_1774; // @[Rob.scala 286:30 Rob.scala 286:30]
  wire  _GEN_1831 = 3'h7 == io_wb_info_i_1_bits_rob_idx ? 1'h0 : _GEN_1775; // @[Rob.scala 286:30 Rob.scala 286:30]
  wire  _GEN_1832 = 3'h0 == io_wb_info_i_1_bits_rob_idx ? 1'h0 : _GEN_1776; // @[Rob.scala 287:34 Rob.scala 287:34]
  wire  _GEN_1833 = 3'h1 == io_wb_info_i_1_bits_rob_idx ? 1'h0 : _GEN_1777; // @[Rob.scala 287:34 Rob.scala 287:34]
  wire  _GEN_1834 = 3'h2 == io_wb_info_i_1_bits_rob_idx ? 1'h0 : _GEN_1778; // @[Rob.scala 287:34 Rob.scala 287:34]
  wire  _GEN_1835 = 3'h3 == io_wb_info_i_1_bits_rob_idx ? 1'h0 : _GEN_1779; // @[Rob.scala 287:34 Rob.scala 287:34]
  wire  _GEN_1836 = 3'h4 == io_wb_info_i_1_bits_rob_idx ? 1'h0 : _GEN_1780; // @[Rob.scala 287:34 Rob.scala 287:34]
  wire  _GEN_1837 = 3'h5 == io_wb_info_i_1_bits_rob_idx ? 1'h0 : _GEN_1781; // @[Rob.scala 287:34 Rob.scala 287:34]
  wire  _GEN_1838 = 3'h6 == io_wb_info_i_1_bits_rob_idx ? 1'h0 : _GEN_1782; // @[Rob.scala 287:34 Rob.scala 287:34]
  wire  _GEN_1839 = 3'h7 == io_wb_info_i_1_bits_rob_idx ? 1'h0 : _GEN_1783; // @[Rob.scala 287:34 Rob.scala 287:34]
  wire  _GEN_1840 = 3'h0 == io_wb_info_i_1_bits_rob_idx ? 1'h0 : _GEN_1784; // @[Rob.scala 288:38 Rob.scala 288:38]
  wire  _GEN_1841 = 3'h1 == io_wb_info_i_1_bits_rob_idx ? 1'h0 : _GEN_1785; // @[Rob.scala 288:38 Rob.scala 288:38]
  wire  _GEN_1842 = 3'h2 == io_wb_info_i_1_bits_rob_idx ? 1'h0 : _GEN_1786; // @[Rob.scala 288:38 Rob.scala 288:38]
  wire  _GEN_1843 = 3'h3 == io_wb_info_i_1_bits_rob_idx ? 1'h0 : _GEN_1787; // @[Rob.scala 288:38 Rob.scala 288:38]
  wire  _GEN_1844 = 3'h4 == io_wb_info_i_1_bits_rob_idx ? 1'h0 : _GEN_1788; // @[Rob.scala 288:38 Rob.scala 288:38]
  wire  _GEN_1845 = 3'h5 == io_wb_info_i_1_bits_rob_idx ? 1'h0 : _GEN_1789; // @[Rob.scala 288:38 Rob.scala 288:38]
  wire  _GEN_1846 = 3'h6 == io_wb_info_i_1_bits_rob_idx ? 1'h0 : _GEN_1790; // @[Rob.scala 288:38 Rob.scala 288:38]
  wire  _GEN_1847 = 3'h7 == io_wb_info_i_1_bits_rob_idx ? 1'h0 : _GEN_1791; // @[Rob.scala 288:38 Rob.scala 288:38]
  wire [31:0] _GEN_1848 = 3'h0 == io_wb_info_i_1_bits_rob_idx ? 32'h0 : _GEN_1792; // @[Rob.scala 289:34 Rob.scala 289:34]
  wire [31:0] _GEN_1849 = 3'h1 == io_wb_info_i_1_bits_rob_idx ? 32'h0 : _GEN_1793; // @[Rob.scala 289:34 Rob.scala 289:34]
  wire [31:0] _GEN_1850 = 3'h2 == io_wb_info_i_1_bits_rob_idx ? 32'h0 : _GEN_1794; // @[Rob.scala 289:34 Rob.scala 289:34]
  wire [31:0] _GEN_1851 = 3'h3 == io_wb_info_i_1_bits_rob_idx ? 32'h0 : _GEN_1795; // @[Rob.scala 289:34 Rob.scala 289:34]
  wire [31:0] _GEN_1852 = 3'h4 == io_wb_info_i_1_bits_rob_idx ? 32'h0 : _GEN_1796; // @[Rob.scala 289:34 Rob.scala 289:34]
  wire [31:0] _GEN_1853 = 3'h5 == io_wb_info_i_1_bits_rob_idx ? 32'h0 : _GEN_1797; // @[Rob.scala 289:34 Rob.scala 289:34]
  wire [31:0] _GEN_1854 = 3'h6 == io_wb_info_i_1_bits_rob_idx ? 32'h0 : _GEN_1798; // @[Rob.scala 289:34 Rob.scala 289:34]
  wire [31:0] _GEN_1855 = 3'h7 == io_wb_info_i_1_bits_rob_idx ? 32'h0 : _GEN_1799; // @[Rob.scala 289:34 Rob.scala 289:34]
  wire [31:0] _GEN_1856 = io_wb_info_i_1_valid & _GEN_1807 & _T_21 ? _GEN_1808 : _GEN_1752; // @[Rob.scala 283:75]
  wire [31:0] _GEN_1857 = io_wb_info_i_1_valid & _GEN_1807 & _T_21 ? _GEN_1809 : _GEN_1753; // @[Rob.scala 283:75]
  wire [31:0] _GEN_1858 = io_wb_info_i_1_valid & _GEN_1807 & _T_21 ? _GEN_1810 : _GEN_1754; // @[Rob.scala 283:75]
  wire [31:0] _GEN_1859 = io_wb_info_i_1_valid & _GEN_1807 & _T_21 ? _GEN_1811 : _GEN_1755; // @[Rob.scala 283:75]
  wire [31:0] _GEN_1860 = io_wb_info_i_1_valid & _GEN_1807 & _T_21 ? _GEN_1812 : _GEN_1756; // @[Rob.scala 283:75]
  wire [31:0] _GEN_1861 = io_wb_info_i_1_valid & _GEN_1807 & _T_21 ? _GEN_1813 : _GEN_1757; // @[Rob.scala 283:75]
  wire [31:0] _GEN_1862 = io_wb_info_i_1_valid & _GEN_1807 & _T_21 ? _GEN_1814 : _GEN_1758; // @[Rob.scala 283:75]
  wire [31:0] _GEN_1863 = io_wb_info_i_1_valid & _GEN_1807 & _T_21 ? _GEN_1815 : _GEN_1759; // @[Rob.scala 283:75]
  wire  _GEN_1864 = io_wb_info_i_1_valid & _GEN_1807 & _T_21 ? _GEN_1816 : _GEN_1760; // @[Rob.scala 283:75]
  wire  _GEN_1865 = io_wb_info_i_1_valid & _GEN_1807 & _T_21 ? _GEN_1817 : _GEN_1761; // @[Rob.scala 283:75]
  wire  _GEN_1866 = io_wb_info_i_1_valid & _GEN_1807 & _T_21 ? _GEN_1818 : _GEN_1762; // @[Rob.scala 283:75]
  wire  _GEN_1867 = io_wb_info_i_1_valid & _GEN_1807 & _T_21 ? _GEN_1819 : _GEN_1763; // @[Rob.scala 283:75]
  wire  _GEN_1868 = io_wb_info_i_1_valid & _GEN_1807 & _T_21 ? _GEN_1820 : _GEN_1764; // @[Rob.scala 283:75]
  wire  _GEN_1869 = io_wb_info_i_1_valid & _GEN_1807 & _T_21 ? _GEN_1821 : _GEN_1765; // @[Rob.scala 283:75]
  wire  _GEN_1870 = io_wb_info_i_1_valid & _GEN_1807 & _T_21 ? _GEN_1822 : _GEN_1766; // @[Rob.scala 283:75]
  wire  _GEN_1871 = io_wb_info_i_1_valid & _GEN_1807 & _T_21 ? _GEN_1823 : _GEN_1767; // @[Rob.scala 283:75]
  wire  _GEN_1872 = io_wb_info_i_1_valid & _GEN_1807 & _T_21 ? _GEN_1824 : _GEN_1768; // @[Rob.scala 283:75]
  wire  _GEN_1873 = io_wb_info_i_1_valid & _GEN_1807 & _T_21 ? _GEN_1825 : _GEN_1769; // @[Rob.scala 283:75]
  wire  _GEN_1874 = io_wb_info_i_1_valid & _GEN_1807 & _T_21 ? _GEN_1826 : _GEN_1770; // @[Rob.scala 283:75]
  wire  _GEN_1875 = io_wb_info_i_1_valid & _GEN_1807 & _T_21 ? _GEN_1827 : _GEN_1771; // @[Rob.scala 283:75]
  wire  _GEN_1876 = io_wb_info_i_1_valid & _GEN_1807 & _T_21 ? _GEN_1828 : _GEN_1772; // @[Rob.scala 283:75]
  wire  _GEN_1877 = io_wb_info_i_1_valid & _GEN_1807 & _T_21 ? _GEN_1829 : _GEN_1773; // @[Rob.scala 283:75]
  wire  _GEN_1878 = io_wb_info_i_1_valid & _GEN_1807 & _T_21 ? _GEN_1830 : _GEN_1774; // @[Rob.scala 283:75]
  wire  _GEN_1879 = io_wb_info_i_1_valid & _GEN_1807 & _T_21 ? _GEN_1831 : _GEN_1775; // @[Rob.scala 283:75]
  wire  _GEN_1880 = io_wb_info_i_1_valid & _GEN_1807 & _T_21 ? _GEN_1832 : _GEN_1776; // @[Rob.scala 283:75]
  wire  _GEN_1881 = io_wb_info_i_1_valid & _GEN_1807 & _T_21 ? _GEN_1833 : _GEN_1777; // @[Rob.scala 283:75]
  wire  _GEN_1882 = io_wb_info_i_1_valid & _GEN_1807 & _T_21 ? _GEN_1834 : _GEN_1778; // @[Rob.scala 283:75]
  wire  _GEN_1883 = io_wb_info_i_1_valid & _GEN_1807 & _T_21 ? _GEN_1835 : _GEN_1779; // @[Rob.scala 283:75]
  wire  _GEN_1884 = io_wb_info_i_1_valid & _GEN_1807 & _T_21 ? _GEN_1836 : _GEN_1780; // @[Rob.scala 283:75]
  wire  _GEN_1885 = io_wb_info_i_1_valid & _GEN_1807 & _T_21 ? _GEN_1837 : _GEN_1781; // @[Rob.scala 283:75]
  wire  _GEN_1886 = io_wb_info_i_1_valid & _GEN_1807 & _T_21 ? _GEN_1838 : _GEN_1782; // @[Rob.scala 283:75]
  wire  _GEN_1887 = io_wb_info_i_1_valid & _GEN_1807 & _T_21 ? _GEN_1839 : _GEN_1783; // @[Rob.scala 283:75]
  wire  _GEN_1888 = io_wb_info_i_1_valid & _GEN_1807 & _T_21 ? _GEN_1840 : _GEN_1784; // @[Rob.scala 283:75]
  wire  _GEN_1889 = io_wb_info_i_1_valid & _GEN_1807 & _T_21 ? _GEN_1841 : _GEN_1785; // @[Rob.scala 283:75]
  wire  _GEN_1890 = io_wb_info_i_1_valid & _GEN_1807 & _T_21 ? _GEN_1842 : _GEN_1786; // @[Rob.scala 283:75]
  wire  _GEN_1891 = io_wb_info_i_1_valid & _GEN_1807 & _T_21 ? _GEN_1843 : _GEN_1787; // @[Rob.scala 283:75]
  wire  _GEN_1892 = io_wb_info_i_1_valid & _GEN_1807 & _T_21 ? _GEN_1844 : _GEN_1788; // @[Rob.scala 283:75]
  wire  _GEN_1893 = io_wb_info_i_1_valid & _GEN_1807 & _T_21 ? _GEN_1845 : _GEN_1789; // @[Rob.scala 283:75]
  wire  _GEN_1894 = io_wb_info_i_1_valid & _GEN_1807 & _T_21 ? _GEN_1846 : _GEN_1790; // @[Rob.scala 283:75]
  wire  _GEN_1895 = io_wb_info_i_1_valid & _GEN_1807 & _T_21 ? _GEN_1847 : _GEN_1791; // @[Rob.scala 283:75]
  wire [31:0] _GEN_1896 = io_wb_info_i_1_valid & _GEN_1807 & _T_21 ? _GEN_1848 : _GEN_1792; // @[Rob.scala 283:75]
  wire [31:0] _GEN_1897 = io_wb_info_i_1_valid & _GEN_1807 & _T_21 ? _GEN_1849 : _GEN_1793; // @[Rob.scala 283:75]
  wire [31:0] _GEN_1898 = io_wb_info_i_1_valid & _GEN_1807 & _T_21 ? _GEN_1850 : _GEN_1794; // @[Rob.scala 283:75]
  wire [31:0] _GEN_1899 = io_wb_info_i_1_valid & _GEN_1807 & _T_21 ? _GEN_1851 : _GEN_1795; // @[Rob.scala 283:75]
  wire [31:0] _GEN_1900 = io_wb_info_i_1_valid & _GEN_1807 & _T_21 ? _GEN_1852 : _GEN_1796; // @[Rob.scala 283:75]
  wire [31:0] _GEN_1901 = io_wb_info_i_1_valid & _GEN_1807 & _T_21 ? _GEN_1853 : _GEN_1797; // @[Rob.scala 283:75]
  wire [31:0] _GEN_1902 = io_wb_info_i_1_valid & _GEN_1807 & _T_21 ? _GEN_1854 : _GEN_1798; // @[Rob.scala 283:75]
  wire [31:0] _GEN_1903 = io_wb_info_i_1_valid & _GEN_1807 & _T_21 ? _GEN_1855 : _GEN_1799; // @[Rob.scala 283:75]
  wire  _GEN_1905 = 3'h1 == io_wb_info_i_2_bits_rob_idx ? rob_info_1_is_valid : rob_info_0_is_valid; // @[Rob.scala 283:31 Rob.scala 283:31]
  wire  _GEN_1906 = 3'h2 == io_wb_info_i_2_bits_rob_idx ? rob_info_2_is_valid : _GEN_1905; // @[Rob.scala 283:31 Rob.scala 283:31]
  wire  _GEN_1907 = 3'h3 == io_wb_info_i_2_bits_rob_idx ? rob_info_3_is_valid : _GEN_1906; // @[Rob.scala 283:31 Rob.scala 283:31]
  wire  _GEN_1908 = 3'h4 == io_wb_info_i_2_bits_rob_idx ? rob_info_4_is_valid : _GEN_1907; // @[Rob.scala 283:31 Rob.scala 283:31]
  wire  _GEN_1909 = 3'h5 == io_wb_info_i_2_bits_rob_idx ? rob_info_5_is_valid : _GEN_1908; // @[Rob.scala 283:31 Rob.scala 283:31]
  wire  _GEN_1910 = 3'h6 == io_wb_info_i_2_bits_rob_idx ? rob_info_6_is_valid : _GEN_1909; // @[Rob.scala 283:31 Rob.scala 283:31]
  wire  _GEN_1911 = 3'h7 == io_wb_info_i_2_bits_rob_idx ? rob_info_7_is_valid : _GEN_1910; // @[Rob.scala 283:31 Rob.scala 283:31]
  wire [31:0] _GEN_1912 = 3'h0 == io_wb_info_i_2_bits_rob_idx ? io_wb_info_i_2_bits_data : _GEN_1856; // @[Rob.scala 284:37 Rob.scala 284:37]
  wire [31:0] _GEN_1913 = 3'h1 == io_wb_info_i_2_bits_rob_idx ? io_wb_info_i_2_bits_data : _GEN_1857; // @[Rob.scala 284:37 Rob.scala 284:37]
  wire [31:0] _GEN_1914 = 3'h2 == io_wb_info_i_2_bits_rob_idx ? io_wb_info_i_2_bits_data : _GEN_1858; // @[Rob.scala 284:37 Rob.scala 284:37]
  wire [31:0] _GEN_1915 = 3'h3 == io_wb_info_i_2_bits_rob_idx ? io_wb_info_i_2_bits_data : _GEN_1859; // @[Rob.scala 284:37 Rob.scala 284:37]
  wire [31:0] _GEN_1916 = 3'h4 == io_wb_info_i_2_bits_rob_idx ? io_wb_info_i_2_bits_data : _GEN_1860; // @[Rob.scala 284:37 Rob.scala 284:37]
  wire [31:0] _GEN_1917 = 3'h5 == io_wb_info_i_2_bits_rob_idx ? io_wb_info_i_2_bits_data : _GEN_1861; // @[Rob.scala 284:37 Rob.scala 284:37]
  wire [31:0] _GEN_1918 = 3'h6 == io_wb_info_i_2_bits_rob_idx ? io_wb_info_i_2_bits_data : _GEN_1862; // @[Rob.scala 284:37 Rob.scala 284:37]
  wire [31:0] _GEN_1919 = 3'h7 == io_wb_info_i_2_bits_rob_idx ? io_wb_info_i_2_bits_data : _GEN_1863; // @[Rob.scala 284:37 Rob.scala 284:37]
  wire  _GEN_1920 = 3'h0 == io_wb_info_i_2_bits_rob_idx | _GEN_1864; // @[Rob.scala 285:38 Rob.scala 285:38]
  wire  _GEN_1921 = 3'h1 == io_wb_info_i_2_bits_rob_idx | _GEN_1865; // @[Rob.scala 285:38 Rob.scala 285:38]
  wire  _GEN_1922 = 3'h2 == io_wb_info_i_2_bits_rob_idx | _GEN_1866; // @[Rob.scala 285:38 Rob.scala 285:38]
  wire  _GEN_1923 = 3'h3 == io_wb_info_i_2_bits_rob_idx | _GEN_1867; // @[Rob.scala 285:38 Rob.scala 285:38]
  wire  _GEN_1924 = 3'h4 == io_wb_info_i_2_bits_rob_idx | _GEN_1868; // @[Rob.scala 285:38 Rob.scala 285:38]
  wire  _GEN_1925 = 3'h5 == io_wb_info_i_2_bits_rob_idx | _GEN_1869; // @[Rob.scala 285:38 Rob.scala 285:38]
  wire  _GEN_1926 = 3'h6 == io_wb_info_i_2_bits_rob_idx | _GEN_1870; // @[Rob.scala 285:38 Rob.scala 285:38]
  wire  _GEN_1927 = 3'h7 == io_wb_info_i_2_bits_rob_idx | _GEN_1871; // @[Rob.scala 285:38 Rob.scala 285:38]
  wire  _GEN_1928 = 3'h0 == io_wb_info_i_2_bits_rob_idx ? 1'h0 : _GEN_1872; // @[Rob.scala 286:30 Rob.scala 286:30]
  wire  _GEN_1929 = 3'h1 == io_wb_info_i_2_bits_rob_idx ? 1'h0 : _GEN_1873; // @[Rob.scala 286:30 Rob.scala 286:30]
  wire  _GEN_1930 = 3'h2 == io_wb_info_i_2_bits_rob_idx ? 1'h0 : _GEN_1874; // @[Rob.scala 286:30 Rob.scala 286:30]
  wire  _GEN_1931 = 3'h3 == io_wb_info_i_2_bits_rob_idx ? 1'h0 : _GEN_1875; // @[Rob.scala 286:30 Rob.scala 286:30]
  wire  _GEN_1932 = 3'h4 == io_wb_info_i_2_bits_rob_idx ? 1'h0 : _GEN_1876; // @[Rob.scala 286:30 Rob.scala 286:30]
  wire  _GEN_1933 = 3'h5 == io_wb_info_i_2_bits_rob_idx ? 1'h0 : _GEN_1877; // @[Rob.scala 286:30 Rob.scala 286:30]
  wire  _GEN_1934 = 3'h6 == io_wb_info_i_2_bits_rob_idx ? 1'h0 : _GEN_1878; // @[Rob.scala 286:30 Rob.scala 286:30]
  wire  _GEN_1935 = 3'h7 == io_wb_info_i_2_bits_rob_idx ? 1'h0 : _GEN_1879; // @[Rob.scala 286:30 Rob.scala 286:30]
  wire  _GEN_1936 = 3'h0 == io_wb_info_i_2_bits_rob_idx ? io_wb_info_i_2_bits_is_taken : _GEN_1880; // @[Rob.scala 287:34 Rob.scala 287:34]
  wire  _GEN_1937 = 3'h1 == io_wb_info_i_2_bits_rob_idx ? io_wb_info_i_2_bits_is_taken : _GEN_1881; // @[Rob.scala 287:34 Rob.scala 287:34]
  wire  _GEN_1938 = 3'h2 == io_wb_info_i_2_bits_rob_idx ? io_wb_info_i_2_bits_is_taken : _GEN_1882; // @[Rob.scala 287:34 Rob.scala 287:34]
  wire  _GEN_1939 = 3'h3 == io_wb_info_i_2_bits_rob_idx ? io_wb_info_i_2_bits_is_taken : _GEN_1883; // @[Rob.scala 287:34 Rob.scala 287:34]
  wire  _GEN_1940 = 3'h4 == io_wb_info_i_2_bits_rob_idx ? io_wb_info_i_2_bits_is_taken : _GEN_1884; // @[Rob.scala 287:34 Rob.scala 287:34]
  wire  _GEN_1941 = 3'h5 == io_wb_info_i_2_bits_rob_idx ? io_wb_info_i_2_bits_is_taken : _GEN_1885; // @[Rob.scala 287:34 Rob.scala 287:34]
  wire  _GEN_1942 = 3'h6 == io_wb_info_i_2_bits_rob_idx ? io_wb_info_i_2_bits_is_taken : _GEN_1886; // @[Rob.scala 287:34 Rob.scala 287:34]
  wire  _GEN_1943 = 3'h7 == io_wb_info_i_2_bits_rob_idx ? io_wb_info_i_2_bits_is_taken : _GEN_1887; // @[Rob.scala 287:34 Rob.scala 287:34]
  wire  _GEN_1944 = 3'h0 == io_wb_info_i_2_bits_rob_idx ? io_wb_info_i_2_bits_predict_miss : _GEN_1888; // @[Rob.scala 288:38 Rob.scala 288:38]
  wire  _GEN_1945 = 3'h1 == io_wb_info_i_2_bits_rob_idx ? io_wb_info_i_2_bits_predict_miss : _GEN_1889; // @[Rob.scala 288:38 Rob.scala 288:38]
  wire  _GEN_1946 = 3'h2 == io_wb_info_i_2_bits_rob_idx ? io_wb_info_i_2_bits_predict_miss : _GEN_1890; // @[Rob.scala 288:38 Rob.scala 288:38]
  wire  _GEN_1947 = 3'h3 == io_wb_info_i_2_bits_rob_idx ? io_wb_info_i_2_bits_predict_miss : _GEN_1891; // @[Rob.scala 288:38 Rob.scala 288:38]
  wire  _GEN_1948 = 3'h4 == io_wb_info_i_2_bits_rob_idx ? io_wb_info_i_2_bits_predict_miss : _GEN_1892; // @[Rob.scala 288:38 Rob.scala 288:38]
  wire  _GEN_1949 = 3'h5 == io_wb_info_i_2_bits_rob_idx ? io_wb_info_i_2_bits_predict_miss : _GEN_1893; // @[Rob.scala 288:38 Rob.scala 288:38]
  wire  _GEN_1950 = 3'h6 == io_wb_info_i_2_bits_rob_idx ? io_wb_info_i_2_bits_predict_miss : _GEN_1894; // @[Rob.scala 288:38 Rob.scala 288:38]
  wire  _GEN_1951 = 3'h7 == io_wb_info_i_2_bits_rob_idx ? io_wb_info_i_2_bits_predict_miss : _GEN_1895; // @[Rob.scala 288:38 Rob.scala 288:38]
  wire [31:0] _GEN_1952 = 3'h0 == io_wb_info_i_2_bits_rob_idx ? io_wb_info_i_2_bits_target_addr : _GEN_1896; // @[Rob.scala 289:34 Rob.scala 289:34]
  wire [31:0] _GEN_1953 = 3'h1 == io_wb_info_i_2_bits_rob_idx ? io_wb_info_i_2_bits_target_addr : _GEN_1897; // @[Rob.scala 289:34 Rob.scala 289:34]
  wire [31:0] _GEN_1954 = 3'h2 == io_wb_info_i_2_bits_rob_idx ? io_wb_info_i_2_bits_target_addr : _GEN_1898; // @[Rob.scala 289:34 Rob.scala 289:34]
  wire [31:0] _GEN_1955 = 3'h3 == io_wb_info_i_2_bits_rob_idx ? io_wb_info_i_2_bits_target_addr : _GEN_1899; // @[Rob.scala 289:34 Rob.scala 289:34]
  wire [31:0] _GEN_1956 = 3'h4 == io_wb_info_i_2_bits_rob_idx ? io_wb_info_i_2_bits_target_addr : _GEN_1900; // @[Rob.scala 289:34 Rob.scala 289:34]
  wire [31:0] _GEN_1957 = 3'h5 == io_wb_info_i_2_bits_rob_idx ? io_wb_info_i_2_bits_target_addr : _GEN_1901; // @[Rob.scala 289:34 Rob.scala 289:34]
  wire [31:0] _GEN_1958 = 3'h6 == io_wb_info_i_2_bits_rob_idx ? io_wb_info_i_2_bits_target_addr : _GEN_1902; // @[Rob.scala 289:34 Rob.scala 289:34]
  wire [31:0] _GEN_1959 = 3'h7 == io_wb_info_i_2_bits_rob_idx ? io_wb_info_i_2_bits_target_addr : _GEN_1903; // @[Rob.scala 289:34 Rob.scala 289:34]
  wire [31:0] _GEN_1960 = io_wb_info_i_2_valid & _GEN_1911 & _T_21 ? _GEN_1912 : _GEN_1856; // @[Rob.scala 283:75]
  wire [31:0] _GEN_1961 = io_wb_info_i_2_valid & _GEN_1911 & _T_21 ? _GEN_1913 : _GEN_1857; // @[Rob.scala 283:75]
  wire [31:0] _GEN_1962 = io_wb_info_i_2_valid & _GEN_1911 & _T_21 ? _GEN_1914 : _GEN_1858; // @[Rob.scala 283:75]
  wire [31:0] _GEN_1963 = io_wb_info_i_2_valid & _GEN_1911 & _T_21 ? _GEN_1915 : _GEN_1859; // @[Rob.scala 283:75]
  wire [31:0] _GEN_1964 = io_wb_info_i_2_valid & _GEN_1911 & _T_21 ? _GEN_1916 : _GEN_1860; // @[Rob.scala 283:75]
  wire [31:0] _GEN_1965 = io_wb_info_i_2_valid & _GEN_1911 & _T_21 ? _GEN_1917 : _GEN_1861; // @[Rob.scala 283:75]
  wire [31:0] _GEN_1966 = io_wb_info_i_2_valid & _GEN_1911 & _T_21 ? _GEN_1918 : _GEN_1862; // @[Rob.scala 283:75]
  wire [31:0] _GEN_1967 = io_wb_info_i_2_valid & _GEN_1911 & _T_21 ? _GEN_1919 : _GEN_1863; // @[Rob.scala 283:75]
  wire  _GEN_1968 = io_wb_info_i_2_valid & _GEN_1911 & _T_21 ? _GEN_1920 : _GEN_1864; // @[Rob.scala 283:75]
  wire  _GEN_1969 = io_wb_info_i_2_valid & _GEN_1911 & _T_21 ? _GEN_1921 : _GEN_1865; // @[Rob.scala 283:75]
  wire  _GEN_1970 = io_wb_info_i_2_valid & _GEN_1911 & _T_21 ? _GEN_1922 : _GEN_1866; // @[Rob.scala 283:75]
  wire  _GEN_1971 = io_wb_info_i_2_valid & _GEN_1911 & _T_21 ? _GEN_1923 : _GEN_1867; // @[Rob.scala 283:75]
  wire  _GEN_1972 = io_wb_info_i_2_valid & _GEN_1911 & _T_21 ? _GEN_1924 : _GEN_1868; // @[Rob.scala 283:75]
  wire  _GEN_1973 = io_wb_info_i_2_valid & _GEN_1911 & _T_21 ? _GEN_1925 : _GEN_1869; // @[Rob.scala 283:75]
  wire  _GEN_1974 = io_wb_info_i_2_valid & _GEN_1911 & _T_21 ? _GEN_1926 : _GEN_1870; // @[Rob.scala 283:75]
  wire  _GEN_1975 = io_wb_info_i_2_valid & _GEN_1911 & _T_21 ? _GEN_1927 : _GEN_1871; // @[Rob.scala 283:75]
  wire  _GEN_1976 = io_wb_info_i_2_valid & _GEN_1911 & _T_21 ? _GEN_1928 : _GEN_1872; // @[Rob.scala 283:75]
  wire  _GEN_1977 = io_wb_info_i_2_valid & _GEN_1911 & _T_21 ? _GEN_1929 : _GEN_1873; // @[Rob.scala 283:75]
  wire  _GEN_1978 = io_wb_info_i_2_valid & _GEN_1911 & _T_21 ? _GEN_1930 : _GEN_1874; // @[Rob.scala 283:75]
  wire  _GEN_1979 = io_wb_info_i_2_valid & _GEN_1911 & _T_21 ? _GEN_1931 : _GEN_1875; // @[Rob.scala 283:75]
  wire  _GEN_1980 = io_wb_info_i_2_valid & _GEN_1911 & _T_21 ? _GEN_1932 : _GEN_1876; // @[Rob.scala 283:75]
  wire  _GEN_1981 = io_wb_info_i_2_valid & _GEN_1911 & _T_21 ? _GEN_1933 : _GEN_1877; // @[Rob.scala 283:75]
  wire  _GEN_1982 = io_wb_info_i_2_valid & _GEN_1911 & _T_21 ? _GEN_1934 : _GEN_1878; // @[Rob.scala 283:75]
  wire  _GEN_1983 = io_wb_info_i_2_valid & _GEN_1911 & _T_21 ? _GEN_1935 : _GEN_1879; // @[Rob.scala 283:75]
  wire  _GEN_1984 = io_wb_info_i_2_valid & _GEN_1911 & _T_21 ? _GEN_1936 : _GEN_1880; // @[Rob.scala 283:75]
  wire  _GEN_1985 = io_wb_info_i_2_valid & _GEN_1911 & _T_21 ? _GEN_1937 : _GEN_1881; // @[Rob.scala 283:75]
  wire  _GEN_1986 = io_wb_info_i_2_valid & _GEN_1911 & _T_21 ? _GEN_1938 : _GEN_1882; // @[Rob.scala 283:75]
  wire  _GEN_1987 = io_wb_info_i_2_valid & _GEN_1911 & _T_21 ? _GEN_1939 : _GEN_1883; // @[Rob.scala 283:75]
  wire  _GEN_1988 = io_wb_info_i_2_valid & _GEN_1911 & _T_21 ? _GEN_1940 : _GEN_1884; // @[Rob.scala 283:75]
  wire  _GEN_1989 = io_wb_info_i_2_valid & _GEN_1911 & _T_21 ? _GEN_1941 : _GEN_1885; // @[Rob.scala 283:75]
  wire  _GEN_1990 = io_wb_info_i_2_valid & _GEN_1911 & _T_21 ? _GEN_1942 : _GEN_1886; // @[Rob.scala 283:75]
  wire  _GEN_1991 = io_wb_info_i_2_valid & _GEN_1911 & _T_21 ? _GEN_1943 : _GEN_1887; // @[Rob.scala 283:75]
  wire  _GEN_1992 = io_wb_info_i_2_valid & _GEN_1911 & _T_21 ? _GEN_1944 : _GEN_1888; // @[Rob.scala 283:75]
  wire  _GEN_1993 = io_wb_info_i_2_valid & _GEN_1911 & _T_21 ? _GEN_1945 : _GEN_1889; // @[Rob.scala 283:75]
  wire  _GEN_1994 = io_wb_info_i_2_valid & _GEN_1911 & _T_21 ? _GEN_1946 : _GEN_1890; // @[Rob.scala 283:75]
  wire  _GEN_1995 = io_wb_info_i_2_valid & _GEN_1911 & _T_21 ? _GEN_1947 : _GEN_1891; // @[Rob.scala 283:75]
  wire  _GEN_1996 = io_wb_info_i_2_valid & _GEN_1911 & _T_21 ? _GEN_1948 : _GEN_1892; // @[Rob.scala 283:75]
  wire  _GEN_1997 = io_wb_info_i_2_valid & _GEN_1911 & _T_21 ? _GEN_1949 : _GEN_1893; // @[Rob.scala 283:75]
  wire  _GEN_1998 = io_wb_info_i_2_valid & _GEN_1911 & _T_21 ? _GEN_1950 : _GEN_1894; // @[Rob.scala 283:75]
  wire  _GEN_1999 = io_wb_info_i_2_valid & _GEN_1911 & _T_21 ? _GEN_1951 : _GEN_1895; // @[Rob.scala 283:75]
  wire [31:0] _GEN_2000 = io_wb_info_i_2_valid & _GEN_1911 & _T_21 ? _GEN_1952 : _GEN_1896; // @[Rob.scala 283:75]
  wire [31:0] _GEN_2001 = io_wb_info_i_2_valid & _GEN_1911 & _T_21 ? _GEN_1953 : _GEN_1897; // @[Rob.scala 283:75]
  wire [31:0] _GEN_2002 = io_wb_info_i_2_valid & _GEN_1911 & _T_21 ? _GEN_1954 : _GEN_1898; // @[Rob.scala 283:75]
  wire [31:0] _GEN_2003 = io_wb_info_i_2_valid & _GEN_1911 & _T_21 ? _GEN_1955 : _GEN_1899; // @[Rob.scala 283:75]
  wire [31:0] _GEN_2004 = io_wb_info_i_2_valid & _GEN_1911 & _T_21 ? _GEN_1956 : _GEN_1900; // @[Rob.scala 283:75]
  wire [31:0] _GEN_2005 = io_wb_info_i_2_valid & _GEN_1911 & _T_21 ? _GEN_1957 : _GEN_1901; // @[Rob.scala 283:75]
  wire [31:0] _GEN_2006 = io_wb_info_i_2_valid & _GEN_1911 & _T_21 ? _GEN_1958 : _GEN_1902; // @[Rob.scala 283:75]
  wire [31:0] _GEN_2007 = io_wb_info_i_2_valid & _GEN_1911 & _T_21 ? _GEN_1959 : _GEN_1903; // @[Rob.scala 283:75]
  wire  _GEN_2009 = 3'h1 == io_wb_info_i_3_bits_rob_idx ? rob_info_1_is_valid : rob_info_0_is_valid; // @[Rob.scala 283:31 Rob.scala 283:31]
  wire  _GEN_2010 = 3'h2 == io_wb_info_i_3_bits_rob_idx ? rob_info_2_is_valid : _GEN_2009; // @[Rob.scala 283:31 Rob.scala 283:31]
  wire  _GEN_2011 = 3'h3 == io_wb_info_i_3_bits_rob_idx ? rob_info_3_is_valid : _GEN_2010; // @[Rob.scala 283:31 Rob.scala 283:31]
  wire  _GEN_2012 = 3'h4 == io_wb_info_i_3_bits_rob_idx ? rob_info_4_is_valid : _GEN_2011; // @[Rob.scala 283:31 Rob.scala 283:31]
  wire  _GEN_2013 = 3'h5 == io_wb_info_i_3_bits_rob_idx ? rob_info_5_is_valid : _GEN_2012; // @[Rob.scala 283:31 Rob.scala 283:31]
  wire  _GEN_2014 = 3'h6 == io_wb_info_i_3_bits_rob_idx ? rob_info_6_is_valid : _GEN_2013; // @[Rob.scala 283:31 Rob.scala 283:31]
  wire  _GEN_2015 = 3'h7 == io_wb_info_i_3_bits_rob_idx ? rob_info_7_is_valid : _GEN_2014; // @[Rob.scala 283:31 Rob.scala 283:31]
  wire [31:0] _GEN_2016 = 3'h0 == io_wb_info_i_3_bits_rob_idx ? io_wb_info_i_3_bits_data : _GEN_1960; // @[Rob.scala 284:37 Rob.scala 284:37]
  wire [31:0] _GEN_2017 = 3'h1 == io_wb_info_i_3_bits_rob_idx ? io_wb_info_i_3_bits_data : _GEN_1961; // @[Rob.scala 284:37 Rob.scala 284:37]
  wire [31:0] _GEN_2018 = 3'h2 == io_wb_info_i_3_bits_rob_idx ? io_wb_info_i_3_bits_data : _GEN_1962; // @[Rob.scala 284:37 Rob.scala 284:37]
  wire [31:0] _GEN_2019 = 3'h3 == io_wb_info_i_3_bits_rob_idx ? io_wb_info_i_3_bits_data : _GEN_1963; // @[Rob.scala 284:37 Rob.scala 284:37]
  wire [31:0] _GEN_2020 = 3'h4 == io_wb_info_i_3_bits_rob_idx ? io_wb_info_i_3_bits_data : _GEN_1964; // @[Rob.scala 284:37 Rob.scala 284:37]
  wire [31:0] _GEN_2021 = 3'h5 == io_wb_info_i_3_bits_rob_idx ? io_wb_info_i_3_bits_data : _GEN_1965; // @[Rob.scala 284:37 Rob.scala 284:37]
  wire [31:0] _GEN_2022 = 3'h6 == io_wb_info_i_3_bits_rob_idx ? io_wb_info_i_3_bits_data : _GEN_1966; // @[Rob.scala 284:37 Rob.scala 284:37]
  wire [31:0] _GEN_2023 = 3'h7 == io_wb_info_i_3_bits_rob_idx ? io_wb_info_i_3_bits_data : _GEN_1967; // @[Rob.scala 284:37 Rob.scala 284:37]
  wire  _GEN_2024 = 3'h0 == io_wb_info_i_3_bits_rob_idx | _GEN_1968; // @[Rob.scala 285:38 Rob.scala 285:38]
  wire  _GEN_2025 = 3'h1 == io_wb_info_i_3_bits_rob_idx | _GEN_1969; // @[Rob.scala 285:38 Rob.scala 285:38]
  wire  _GEN_2026 = 3'h2 == io_wb_info_i_3_bits_rob_idx | _GEN_1970; // @[Rob.scala 285:38 Rob.scala 285:38]
  wire  _GEN_2027 = 3'h3 == io_wb_info_i_3_bits_rob_idx | _GEN_1971; // @[Rob.scala 285:38 Rob.scala 285:38]
  wire  _GEN_2028 = 3'h4 == io_wb_info_i_3_bits_rob_idx | _GEN_1972; // @[Rob.scala 285:38 Rob.scala 285:38]
  wire  _GEN_2029 = 3'h5 == io_wb_info_i_3_bits_rob_idx | _GEN_1973; // @[Rob.scala 285:38 Rob.scala 285:38]
  wire  _GEN_2030 = 3'h6 == io_wb_info_i_3_bits_rob_idx | _GEN_1974; // @[Rob.scala 285:38 Rob.scala 285:38]
  wire  _GEN_2031 = 3'h7 == io_wb_info_i_3_bits_rob_idx | _GEN_1975; // @[Rob.scala 285:38 Rob.scala 285:38]
  wire  _GEN_2032 = 3'h0 == io_wb_info_i_3_bits_rob_idx ? 1'h0 : _GEN_1976; // @[Rob.scala 286:30 Rob.scala 286:30]
  wire  _GEN_2033 = 3'h1 == io_wb_info_i_3_bits_rob_idx ? 1'h0 : _GEN_1977; // @[Rob.scala 286:30 Rob.scala 286:30]
  wire  _GEN_2034 = 3'h2 == io_wb_info_i_3_bits_rob_idx ? 1'h0 : _GEN_1978; // @[Rob.scala 286:30 Rob.scala 286:30]
  wire  _GEN_2035 = 3'h3 == io_wb_info_i_3_bits_rob_idx ? 1'h0 : _GEN_1979; // @[Rob.scala 286:30 Rob.scala 286:30]
  wire  _GEN_2036 = 3'h4 == io_wb_info_i_3_bits_rob_idx ? 1'h0 : _GEN_1980; // @[Rob.scala 286:30 Rob.scala 286:30]
  wire  _GEN_2037 = 3'h5 == io_wb_info_i_3_bits_rob_idx ? 1'h0 : _GEN_1981; // @[Rob.scala 286:30 Rob.scala 286:30]
  wire  _GEN_2038 = 3'h6 == io_wb_info_i_3_bits_rob_idx ? 1'h0 : _GEN_1982; // @[Rob.scala 286:30 Rob.scala 286:30]
  wire  _GEN_2039 = 3'h7 == io_wb_info_i_3_bits_rob_idx ? 1'h0 : _GEN_1983; // @[Rob.scala 286:30 Rob.scala 286:30]
  wire  _GEN_2040 = 3'h0 == io_wb_info_i_3_bits_rob_idx ? 1'h0 : _GEN_1984; // @[Rob.scala 287:34 Rob.scala 287:34]
  wire  _GEN_2041 = 3'h1 == io_wb_info_i_3_bits_rob_idx ? 1'h0 : _GEN_1985; // @[Rob.scala 287:34 Rob.scala 287:34]
  wire  _GEN_2042 = 3'h2 == io_wb_info_i_3_bits_rob_idx ? 1'h0 : _GEN_1986; // @[Rob.scala 287:34 Rob.scala 287:34]
  wire  _GEN_2043 = 3'h3 == io_wb_info_i_3_bits_rob_idx ? 1'h0 : _GEN_1987; // @[Rob.scala 287:34 Rob.scala 287:34]
  wire  _GEN_2044 = 3'h4 == io_wb_info_i_3_bits_rob_idx ? 1'h0 : _GEN_1988; // @[Rob.scala 287:34 Rob.scala 287:34]
  wire  _GEN_2045 = 3'h5 == io_wb_info_i_3_bits_rob_idx ? 1'h0 : _GEN_1989; // @[Rob.scala 287:34 Rob.scala 287:34]
  wire  _GEN_2046 = 3'h6 == io_wb_info_i_3_bits_rob_idx ? 1'h0 : _GEN_1990; // @[Rob.scala 287:34 Rob.scala 287:34]
  wire  _GEN_2047 = 3'h7 == io_wb_info_i_3_bits_rob_idx ? 1'h0 : _GEN_1991; // @[Rob.scala 287:34 Rob.scala 287:34]
  wire  _GEN_2048 = 3'h0 == io_wb_info_i_3_bits_rob_idx ? 1'h0 : _GEN_1992; // @[Rob.scala 288:38 Rob.scala 288:38]
  wire  _GEN_2049 = 3'h1 == io_wb_info_i_3_bits_rob_idx ? 1'h0 : _GEN_1993; // @[Rob.scala 288:38 Rob.scala 288:38]
  wire  _GEN_2050 = 3'h2 == io_wb_info_i_3_bits_rob_idx ? 1'h0 : _GEN_1994; // @[Rob.scala 288:38 Rob.scala 288:38]
  wire  _GEN_2051 = 3'h3 == io_wb_info_i_3_bits_rob_idx ? 1'h0 : _GEN_1995; // @[Rob.scala 288:38 Rob.scala 288:38]
  wire  _GEN_2052 = 3'h4 == io_wb_info_i_3_bits_rob_idx ? 1'h0 : _GEN_1996; // @[Rob.scala 288:38 Rob.scala 288:38]
  wire  _GEN_2053 = 3'h5 == io_wb_info_i_3_bits_rob_idx ? 1'h0 : _GEN_1997; // @[Rob.scala 288:38 Rob.scala 288:38]
  wire  _GEN_2054 = 3'h6 == io_wb_info_i_3_bits_rob_idx ? 1'h0 : _GEN_1998; // @[Rob.scala 288:38 Rob.scala 288:38]
  wire  _GEN_2055 = 3'h7 == io_wb_info_i_3_bits_rob_idx ? 1'h0 : _GEN_1999; // @[Rob.scala 288:38 Rob.scala 288:38]
  wire [31:0] _GEN_2056 = 3'h0 == io_wb_info_i_3_bits_rob_idx ? 32'h0 : _GEN_2000; // @[Rob.scala 289:34 Rob.scala 289:34]
  wire [31:0] _GEN_2057 = 3'h1 == io_wb_info_i_3_bits_rob_idx ? 32'h0 : _GEN_2001; // @[Rob.scala 289:34 Rob.scala 289:34]
  wire [31:0] _GEN_2058 = 3'h2 == io_wb_info_i_3_bits_rob_idx ? 32'h0 : _GEN_2002; // @[Rob.scala 289:34 Rob.scala 289:34]
  wire [31:0] _GEN_2059 = 3'h3 == io_wb_info_i_3_bits_rob_idx ? 32'h0 : _GEN_2003; // @[Rob.scala 289:34 Rob.scala 289:34]
  wire [31:0] _GEN_2060 = 3'h4 == io_wb_info_i_3_bits_rob_idx ? 32'h0 : _GEN_2004; // @[Rob.scala 289:34 Rob.scala 289:34]
  wire [31:0] _GEN_2061 = 3'h5 == io_wb_info_i_3_bits_rob_idx ? 32'h0 : _GEN_2005; // @[Rob.scala 289:34 Rob.scala 289:34]
  wire [31:0] _GEN_2062 = 3'h6 == io_wb_info_i_3_bits_rob_idx ? 32'h0 : _GEN_2006; // @[Rob.scala 289:34 Rob.scala 289:34]
  wire [31:0] _GEN_2063 = 3'h7 == io_wb_info_i_3_bits_rob_idx ? 32'h0 : _GEN_2007; // @[Rob.scala 289:34 Rob.scala 289:34]
  wire [31:0] _GEN_2064 = io_wb_info_i_3_valid & _GEN_2015 & _T_21 ? _GEN_2016 : _GEN_1960; // @[Rob.scala 283:75]
  wire [31:0] _GEN_2065 = io_wb_info_i_3_valid & _GEN_2015 & _T_21 ? _GEN_2017 : _GEN_1961; // @[Rob.scala 283:75]
  wire [31:0] _GEN_2066 = io_wb_info_i_3_valid & _GEN_2015 & _T_21 ? _GEN_2018 : _GEN_1962; // @[Rob.scala 283:75]
  wire [31:0] _GEN_2067 = io_wb_info_i_3_valid & _GEN_2015 & _T_21 ? _GEN_2019 : _GEN_1963; // @[Rob.scala 283:75]
  wire [31:0] _GEN_2068 = io_wb_info_i_3_valid & _GEN_2015 & _T_21 ? _GEN_2020 : _GEN_1964; // @[Rob.scala 283:75]
  wire [31:0] _GEN_2069 = io_wb_info_i_3_valid & _GEN_2015 & _T_21 ? _GEN_2021 : _GEN_1965; // @[Rob.scala 283:75]
  wire [31:0] _GEN_2070 = io_wb_info_i_3_valid & _GEN_2015 & _T_21 ? _GEN_2022 : _GEN_1966; // @[Rob.scala 283:75]
  wire [31:0] _GEN_2071 = io_wb_info_i_3_valid & _GEN_2015 & _T_21 ? _GEN_2023 : _GEN_1967; // @[Rob.scala 283:75]
  wire  _GEN_2072 = io_wb_info_i_3_valid & _GEN_2015 & _T_21 ? _GEN_2024 : _GEN_1968; // @[Rob.scala 283:75]
  wire  _GEN_2073 = io_wb_info_i_3_valid & _GEN_2015 & _T_21 ? _GEN_2025 : _GEN_1969; // @[Rob.scala 283:75]
  wire  _GEN_2074 = io_wb_info_i_3_valid & _GEN_2015 & _T_21 ? _GEN_2026 : _GEN_1970; // @[Rob.scala 283:75]
  wire  _GEN_2075 = io_wb_info_i_3_valid & _GEN_2015 & _T_21 ? _GEN_2027 : _GEN_1971; // @[Rob.scala 283:75]
  wire  _GEN_2076 = io_wb_info_i_3_valid & _GEN_2015 & _T_21 ? _GEN_2028 : _GEN_1972; // @[Rob.scala 283:75]
  wire  _GEN_2077 = io_wb_info_i_3_valid & _GEN_2015 & _T_21 ? _GEN_2029 : _GEN_1973; // @[Rob.scala 283:75]
  wire  _GEN_2078 = io_wb_info_i_3_valid & _GEN_2015 & _T_21 ? _GEN_2030 : _GEN_1974; // @[Rob.scala 283:75]
  wire  _GEN_2079 = io_wb_info_i_3_valid & _GEN_2015 & _T_21 ? _GEN_2031 : _GEN_1975; // @[Rob.scala 283:75]
  wire  _GEN_2080 = io_wb_info_i_3_valid & _GEN_2015 & _T_21 ? _GEN_2032 : _GEN_1976; // @[Rob.scala 283:75]
  wire  _GEN_2081 = io_wb_info_i_3_valid & _GEN_2015 & _T_21 ? _GEN_2033 : _GEN_1977; // @[Rob.scala 283:75]
  wire  _GEN_2082 = io_wb_info_i_3_valid & _GEN_2015 & _T_21 ? _GEN_2034 : _GEN_1978; // @[Rob.scala 283:75]
  wire  _GEN_2083 = io_wb_info_i_3_valid & _GEN_2015 & _T_21 ? _GEN_2035 : _GEN_1979; // @[Rob.scala 283:75]
  wire  _GEN_2084 = io_wb_info_i_3_valid & _GEN_2015 & _T_21 ? _GEN_2036 : _GEN_1980; // @[Rob.scala 283:75]
  wire  _GEN_2085 = io_wb_info_i_3_valid & _GEN_2015 & _T_21 ? _GEN_2037 : _GEN_1981; // @[Rob.scala 283:75]
  wire  _GEN_2086 = io_wb_info_i_3_valid & _GEN_2015 & _T_21 ? _GEN_2038 : _GEN_1982; // @[Rob.scala 283:75]
  wire  _GEN_2087 = io_wb_info_i_3_valid & _GEN_2015 & _T_21 ? _GEN_2039 : _GEN_1983; // @[Rob.scala 283:75]
  wire  _GEN_2088 = io_wb_info_i_3_valid & _GEN_2015 & _T_21 ? _GEN_2040 : _GEN_1984; // @[Rob.scala 283:75]
  wire  _GEN_2089 = io_wb_info_i_3_valid & _GEN_2015 & _T_21 ? _GEN_2041 : _GEN_1985; // @[Rob.scala 283:75]
  wire  _GEN_2090 = io_wb_info_i_3_valid & _GEN_2015 & _T_21 ? _GEN_2042 : _GEN_1986; // @[Rob.scala 283:75]
  wire  _GEN_2091 = io_wb_info_i_3_valid & _GEN_2015 & _T_21 ? _GEN_2043 : _GEN_1987; // @[Rob.scala 283:75]
  wire  _GEN_2092 = io_wb_info_i_3_valid & _GEN_2015 & _T_21 ? _GEN_2044 : _GEN_1988; // @[Rob.scala 283:75]
  wire  _GEN_2093 = io_wb_info_i_3_valid & _GEN_2015 & _T_21 ? _GEN_2045 : _GEN_1989; // @[Rob.scala 283:75]
  wire  _GEN_2094 = io_wb_info_i_3_valid & _GEN_2015 & _T_21 ? _GEN_2046 : _GEN_1990; // @[Rob.scala 283:75]
  wire  _GEN_2095 = io_wb_info_i_3_valid & _GEN_2015 & _T_21 ? _GEN_2047 : _GEN_1991; // @[Rob.scala 283:75]
  wire  _GEN_2096 = io_wb_info_i_3_valid & _GEN_2015 & _T_21 ? _GEN_2048 : _GEN_1992; // @[Rob.scala 283:75]
  wire  _GEN_2097 = io_wb_info_i_3_valid & _GEN_2015 & _T_21 ? _GEN_2049 : _GEN_1993; // @[Rob.scala 283:75]
  wire  _GEN_2098 = io_wb_info_i_3_valid & _GEN_2015 & _T_21 ? _GEN_2050 : _GEN_1994; // @[Rob.scala 283:75]
  wire  _GEN_2099 = io_wb_info_i_3_valid & _GEN_2015 & _T_21 ? _GEN_2051 : _GEN_1995; // @[Rob.scala 283:75]
  wire  _GEN_2100 = io_wb_info_i_3_valid & _GEN_2015 & _T_21 ? _GEN_2052 : _GEN_1996; // @[Rob.scala 283:75]
  wire  _GEN_2101 = io_wb_info_i_3_valid & _GEN_2015 & _T_21 ? _GEN_2053 : _GEN_1997; // @[Rob.scala 283:75]
  wire  _GEN_2102 = io_wb_info_i_3_valid & _GEN_2015 & _T_21 ? _GEN_2054 : _GEN_1998; // @[Rob.scala 283:75]
  wire  _GEN_2103 = io_wb_info_i_3_valid & _GEN_2015 & _T_21 ? _GEN_2055 : _GEN_1999; // @[Rob.scala 283:75]
  wire [31:0] _GEN_2104 = io_wb_info_i_3_valid & _GEN_2015 & _T_21 ? _GEN_2056 : _GEN_2000; // @[Rob.scala 283:75]
  wire [31:0] _GEN_2105 = io_wb_info_i_3_valid & _GEN_2015 & _T_21 ? _GEN_2057 : _GEN_2001; // @[Rob.scala 283:75]
  wire [31:0] _GEN_2106 = io_wb_info_i_3_valid & _GEN_2015 & _T_21 ? _GEN_2058 : _GEN_2002; // @[Rob.scala 283:75]
  wire [31:0] _GEN_2107 = io_wb_info_i_3_valid & _GEN_2015 & _T_21 ? _GEN_2059 : _GEN_2003; // @[Rob.scala 283:75]
  wire [31:0] _GEN_2108 = io_wb_info_i_3_valid & _GEN_2015 & _T_21 ? _GEN_2060 : _GEN_2004; // @[Rob.scala 283:75]
  wire [31:0] _GEN_2109 = io_wb_info_i_3_valid & _GEN_2015 & _T_21 ? _GEN_2061 : _GEN_2005; // @[Rob.scala 283:75]
  wire [31:0] _GEN_2110 = io_wb_info_i_3_valid & _GEN_2015 & _T_21 ? _GEN_2062 : _GEN_2006; // @[Rob.scala 283:75]
  wire [31:0] _GEN_2111 = io_wb_info_i_3_valid & _GEN_2015 & _T_21 ? _GEN_2063 : _GEN_2007; // @[Rob.scala 283:75]
  wire  _GEN_2113 = 3'h1 == io_wb_info_i_4_bits_rob_idx ? rob_info_1_is_valid : rob_info_0_is_valid; // @[Rob.scala 283:31 Rob.scala 283:31]
  wire  _GEN_2114 = 3'h2 == io_wb_info_i_4_bits_rob_idx ? rob_info_2_is_valid : _GEN_2113; // @[Rob.scala 283:31 Rob.scala 283:31]
  wire  _GEN_2115 = 3'h3 == io_wb_info_i_4_bits_rob_idx ? rob_info_3_is_valid : _GEN_2114; // @[Rob.scala 283:31 Rob.scala 283:31]
  wire  _GEN_2116 = 3'h4 == io_wb_info_i_4_bits_rob_idx ? rob_info_4_is_valid : _GEN_2115; // @[Rob.scala 283:31 Rob.scala 283:31]
  wire  _GEN_2117 = 3'h5 == io_wb_info_i_4_bits_rob_idx ? rob_info_5_is_valid : _GEN_2116; // @[Rob.scala 283:31 Rob.scala 283:31]
  wire  _GEN_2118 = 3'h6 == io_wb_info_i_4_bits_rob_idx ? rob_info_6_is_valid : _GEN_2117; // @[Rob.scala 283:31 Rob.scala 283:31]
  wire  _GEN_2119 = 3'h7 == io_wb_info_i_4_bits_rob_idx ? rob_info_7_is_valid : _GEN_2118; // @[Rob.scala 283:31 Rob.scala 283:31]
  wire [31:0] _GEN_2120 = 3'h0 == io_wb_info_i_4_bits_rob_idx ? io_wb_info_i_4_bits_data : _GEN_2064; // @[Rob.scala 284:37 Rob.scala 284:37]
  wire [31:0] _GEN_2121 = 3'h1 == io_wb_info_i_4_bits_rob_idx ? io_wb_info_i_4_bits_data : _GEN_2065; // @[Rob.scala 284:37 Rob.scala 284:37]
  wire [31:0] _GEN_2122 = 3'h2 == io_wb_info_i_4_bits_rob_idx ? io_wb_info_i_4_bits_data : _GEN_2066; // @[Rob.scala 284:37 Rob.scala 284:37]
  wire [31:0] _GEN_2123 = 3'h3 == io_wb_info_i_4_bits_rob_idx ? io_wb_info_i_4_bits_data : _GEN_2067; // @[Rob.scala 284:37 Rob.scala 284:37]
  wire [31:0] _GEN_2124 = 3'h4 == io_wb_info_i_4_bits_rob_idx ? io_wb_info_i_4_bits_data : _GEN_2068; // @[Rob.scala 284:37 Rob.scala 284:37]
  wire [31:0] _GEN_2125 = 3'h5 == io_wb_info_i_4_bits_rob_idx ? io_wb_info_i_4_bits_data : _GEN_2069; // @[Rob.scala 284:37 Rob.scala 284:37]
  wire [31:0] _GEN_2126 = 3'h6 == io_wb_info_i_4_bits_rob_idx ? io_wb_info_i_4_bits_data : _GEN_2070; // @[Rob.scala 284:37 Rob.scala 284:37]
  wire [31:0] _GEN_2127 = 3'h7 == io_wb_info_i_4_bits_rob_idx ? io_wb_info_i_4_bits_data : _GEN_2071; // @[Rob.scala 284:37 Rob.scala 284:37]
  wire  _GEN_2128 = 3'h0 == io_wb_info_i_4_bits_rob_idx | _GEN_2072; // @[Rob.scala 285:38 Rob.scala 285:38]
  wire  _GEN_2129 = 3'h1 == io_wb_info_i_4_bits_rob_idx | _GEN_2073; // @[Rob.scala 285:38 Rob.scala 285:38]
  wire  _GEN_2130 = 3'h2 == io_wb_info_i_4_bits_rob_idx | _GEN_2074; // @[Rob.scala 285:38 Rob.scala 285:38]
  wire  _GEN_2131 = 3'h3 == io_wb_info_i_4_bits_rob_idx | _GEN_2075; // @[Rob.scala 285:38 Rob.scala 285:38]
  wire  _GEN_2132 = 3'h4 == io_wb_info_i_4_bits_rob_idx | _GEN_2076; // @[Rob.scala 285:38 Rob.scala 285:38]
  wire  _GEN_2133 = 3'h5 == io_wb_info_i_4_bits_rob_idx | _GEN_2077; // @[Rob.scala 285:38 Rob.scala 285:38]
  wire  _GEN_2134 = 3'h6 == io_wb_info_i_4_bits_rob_idx | _GEN_2078; // @[Rob.scala 285:38 Rob.scala 285:38]
  wire  _GEN_2135 = 3'h7 == io_wb_info_i_4_bits_rob_idx | _GEN_2079; // @[Rob.scala 285:38 Rob.scala 285:38]
  wire  _GEN_2136 = 3'h0 == io_wb_info_i_4_bits_rob_idx ? 1'h0 : _GEN_2080; // @[Rob.scala 286:30 Rob.scala 286:30]
  wire  _GEN_2137 = 3'h1 == io_wb_info_i_4_bits_rob_idx ? 1'h0 : _GEN_2081; // @[Rob.scala 286:30 Rob.scala 286:30]
  wire  _GEN_2138 = 3'h2 == io_wb_info_i_4_bits_rob_idx ? 1'h0 : _GEN_2082; // @[Rob.scala 286:30 Rob.scala 286:30]
  wire  _GEN_2139 = 3'h3 == io_wb_info_i_4_bits_rob_idx ? 1'h0 : _GEN_2083; // @[Rob.scala 286:30 Rob.scala 286:30]
  wire  _GEN_2140 = 3'h4 == io_wb_info_i_4_bits_rob_idx ? 1'h0 : _GEN_2084; // @[Rob.scala 286:30 Rob.scala 286:30]
  wire  _GEN_2141 = 3'h5 == io_wb_info_i_4_bits_rob_idx ? 1'h0 : _GEN_2085; // @[Rob.scala 286:30 Rob.scala 286:30]
  wire  _GEN_2142 = 3'h6 == io_wb_info_i_4_bits_rob_idx ? 1'h0 : _GEN_2086; // @[Rob.scala 286:30 Rob.scala 286:30]
  wire  _GEN_2143 = 3'h7 == io_wb_info_i_4_bits_rob_idx ? 1'h0 : _GEN_2087; // @[Rob.scala 286:30 Rob.scala 286:30]
  wire  _GEN_2144 = 3'h0 == io_wb_info_i_4_bits_rob_idx ? 1'h0 : _GEN_2088; // @[Rob.scala 287:34 Rob.scala 287:34]
  wire  _GEN_2145 = 3'h1 == io_wb_info_i_4_bits_rob_idx ? 1'h0 : _GEN_2089; // @[Rob.scala 287:34 Rob.scala 287:34]
  wire  _GEN_2146 = 3'h2 == io_wb_info_i_4_bits_rob_idx ? 1'h0 : _GEN_2090; // @[Rob.scala 287:34 Rob.scala 287:34]
  wire  _GEN_2147 = 3'h3 == io_wb_info_i_4_bits_rob_idx ? 1'h0 : _GEN_2091; // @[Rob.scala 287:34 Rob.scala 287:34]
  wire  _GEN_2148 = 3'h4 == io_wb_info_i_4_bits_rob_idx ? 1'h0 : _GEN_2092; // @[Rob.scala 287:34 Rob.scala 287:34]
  wire  _GEN_2149 = 3'h5 == io_wb_info_i_4_bits_rob_idx ? 1'h0 : _GEN_2093; // @[Rob.scala 287:34 Rob.scala 287:34]
  wire  _GEN_2150 = 3'h6 == io_wb_info_i_4_bits_rob_idx ? 1'h0 : _GEN_2094; // @[Rob.scala 287:34 Rob.scala 287:34]
  wire  _GEN_2151 = 3'h7 == io_wb_info_i_4_bits_rob_idx ? 1'h0 : _GEN_2095; // @[Rob.scala 287:34 Rob.scala 287:34]
  wire  _GEN_2152 = 3'h0 == io_wb_info_i_4_bits_rob_idx ? 1'h0 : _GEN_2096; // @[Rob.scala 288:38 Rob.scala 288:38]
  wire  _GEN_2153 = 3'h1 == io_wb_info_i_4_bits_rob_idx ? 1'h0 : _GEN_2097; // @[Rob.scala 288:38 Rob.scala 288:38]
  wire  _GEN_2154 = 3'h2 == io_wb_info_i_4_bits_rob_idx ? 1'h0 : _GEN_2098; // @[Rob.scala 288:38 Rob.scala 288:38]
  wire  _GEN_2155 = 3'h3 == io_wb_info_i_4_bits_rob_idx ? 1'h0 : _GEN_2099; // @[Rob.scala 288:38 Rob.scala 288:38]
  wire  _GEN_2156 = 3'h4 == io_wb_info_i_4_bits_rob_idx ? 1'h0 : _GEN_2100; // @[Rob.scala 288:38 Rob.scala 288:38]
  wire  _GEN_2157 = 3'h5 == io_wb_info_i_4_bits_rob_idx ? 1'h0 : _GEN_2101; // @[Rob.scala 288:38 Rob.scala 288:38]
  wire  _GEN_2158 = 3'h6 == io_wb_info_i_4_bits_rob_idx ? 1'h0 : _GEN_2102; // @[Rob.scala 288:38 Rob.scala 288:38]
  wire  _GEN_2159 = 3'h7 == io_wb_info_i_4_bits_rob_idx ? 1'h0 : _GEN_2103; // @[Rob.scala 288:38 Rob.scala 288:38]
  wire [31:0] _GEN_2160 = 3'h0 == io_wb_info_i_4_bits_rob_idx ? 32'h0 : _GEN_2104; // @[Rob.scala 289:34 Rob.scala 289:34]
  wire [31:0] _GEN_2161 = 3'h1 == io_wb_info_i_4_bits_rob_idx ? 32'h0 : _GEN_2105; // @[Rob.scala 289:34 Rob.scala 289:34]
  wire [31:0] _GEN_2162 = 3'h2 == io_wb_info_i_4_bits_rob_idx ? 32'h0 : _GEN_2106; // @[Rob.scala 289:34 Rob.scala 289:34]
  wire [31:0] _GEN_2163 = 3'h3 == io_wb_info_i_4_bits_rob_idx ? 32'h0 : _GEN_2107; // @[Rob.scala 289:34 Rob.scala 289:34]
  wire [31:0] _GEN_2164 = 3'h4 == io_wb_info_i_4_bits_rob_idx ? 32'h0 : _GEN_2108; // @[Rob.scala 289:34 Rob.scala 289:34]
  wire [31:0] _GEN_2165 = 3'h5 == io_wb_info_i_4_bits_rob_idx ? 32'h0 : _GEN_2109; // @[Rob.scala 289:34 Rob.scala 289:34]
  wire [31:0] _GEN_2166 = 3'h6 == io_wb_info_i_4_bits_rob_idx ? 32'h0 : _GEN_2110; // @[Rob.scala 289:34 Rob.scala 289:34]
  wire [31:0] _GEN_2167 = 3'h7 == io_wb_info_i_4_bits_rob_idx ? 32'h0 : _GEN_2111; // @[Rob.scala 289:34 Rob.scala 289:34]
  wire [31:0] _GEN_2168 = io_wb_info_i_4_valid & _GEN_2119 & _T_21 ? _GEN_2120 : _GEN_2064; // @[Rob.scala 283:75]
  wire [31:0] _GEN_2169 = io_wb_info_i_4_valid & _GEN_2119 & _T_21 ? _GEN_2121 : _GEN_2065; // @[Rob.scala 283:75]
  wire [31:0] _GEN_2170 = io_wb_info_i_4_valid & _GEN_2119 & _T_21 ? _GEN_2122 : _GEN_2066; // @[Rob.scala 283:75]
  wire [31:0] _GEN_2171 = io_wb_info_i_4_valid & _GEN_2119 & _T_21 ? _GEN_2123 : _GEN_2067; // @[Rob.scala 283:75]
  wire [31:0] _GEN_2172 = io_wb_info_i_4_valid & _GEN_2119 & _T_21 ? _GEN_2124 : _GEN_2068; // @[Rob.scala 283:75]
  wire [31:0] _GEN_2173 = io_wb_info_i_4_valid & _GEN_2119 & _T_21 ? _GEN_2125 : _GEN_2069; // @[Rob.scala 283:75]
  wire [31:0] _GEN_2174 = io_wb_info_i_4_valid & _GEN_2119 & _T_21 ? _GEN_2126 : _GEN_2070; // @[Rob.scala 283:75]
  wire [31:0] _GEN_2175 = io_wb_info_i_4_valid & _GEN_2119 & _T_21 ? _GEN_2127 : _GEN_2071; // @[Rob.scala 283:75]
  wire  _GEN_2176 = io_wb_info_i_4_valid & _GEN_2119 & _T_21 ? _GEN_2128 : _GEN_2072; // @[Rob.scala 283:75]
  wire  _GEN_2177 = io_wb_info_i_4_valid & _GEN_2119 & _T_21 ? _GEN_2129 : _GEN_2073; // @[Rob.scala 283:75]
  wire  _GEN_2178 = io_wb_info_i_4_valid & _GEN_2119 & _T_21 ? _GEN_2130 : _GEN_2074; // @[Rob.scala 283:75]
  wire  _GEN_2179 = io_wb_info_i_4_valid & _GEN_2119 & _T_21 ? _GEN_2131 : _GEN_2075; // @[Rob.scala 283:75]
  wire  _GEN_2180 = io_wb_info_i_4_valid & _GEN_2119 & _T_21 ? _GEN_2132 : _GEN_2076; // @[Rob.scala 283:75]
  wire  _GEN_2181 = io_wb_info_i_4_valid & _GEN_2119 & _T_21 ? _GEN_2133 : _GEN_2077; // @[Rob.scala 283:75]
  wire  _GEN_2182 = io_wb_info_i_4_valid & _GEN_2119 & _T_21 ? _GEN_2134 : _GEN_2078; // @[Rob.scala 283:75]
  wire  _GEN_2183 = io_wb_info_i_4_valid & _GEN_2119 & _T_21 ? _GEN_2135 : _GEN_2079; // @[Rob.scala 283:75]
  wire  _GEN_2184 = io_wb_info_i_4_valid & _GEN_2119 & _T_21 ? _GEN_2136 : _GEN_2080; // @[Rob.scala 283:75]
  wire  _GEN_2185 = io_wb_info_i_4_valid & _GEN_2119 & _T_21 ? _GEN_2137 : _GEN_2081; // @[Rob.scala 283:75]
  wire  _GEN_2186 = io_wb_info_i_4_valid & _GEN_2119 & _T_21 ? _GEN_2138 : _GEN_2082; // @[Rob.scala 283:75]
  wire  _GEN_2187 = io_wb_info_i_4_valid & _GEN_2119 & _T_21 ? _GEN_2139 : _GEN_2083; // @[Rob.scala 283:75]
  wire  _GEN_2188 = io_wb_info_i_4_valid & _GEN_2119 & _T_21 ? _GEN_2140 : _GEN_2084; // @[Rob.scala 283:75]
  wire  _GEN_2189 = io_wb_info_i_4_valid & _GEN_2119 & _T_21 ? _GEN_2141 : _GEN_2085; // @[Rob.scala 283:75]
  wire  _GEN_2190 = io_wb_info_i_4_valid & _GEN_2119 & _T_21 ? _GEN_2142 : _GEN_2086; // @[Rob.scala 283:75]
  wire  _GEN_2191 = io_wb_info_i_4_valid & _GEN_2119 & _T_21 ? _GEN_2143 : _GEN_2087; // @[Rob.scala 283:75]
  wire  _GEN_2192 = io_wb_info_i_4_valid & _GEN_2119 & _T_21 ? _GEN_2144 : _GEN_2088; // @[Rob.scala 283:75]
  wire  _GEN_2193 = io_wb_info_i_4_valid & _GEN_2119 & _T_21 ? _GEN_2145 : _GEN_2089; // @[Rob.scala 283:75]
  wire  _GEN_2194 = io_wb_info_i_4_valid & _GEN_2119 & _T_21 ? _GEN_2146 : _GEN_2090; // @[Rob.scala 283:75]
  wire  _GEN_2195 = io_wb_info_i_4_valid & _GEN_2119 & _T_21 ? _GEN_2147 : _GEN_2091; // @[Rob.scala 283:75]
  wire  _GEN_2196 = io_wb_info_i_4_valid & _GEN_2119 & _T_21 ? _GEN_2148 : _GEN_2092; // @[Rob.scala 283:75]
  wire  _GEN_2197 = io_wb_info_i_4_valid & _GEN_2119 & _T_21 ? _GEN_2149 : _GEN_2093; // @[Rob.scala 283:75]
  wire  _GEN_2198 = io_wb_info_i_4_valid & _GEN_2119 & _T_21 ? _GEN_2150 : _GEN_2094; // @[Rob.scala 283:75]
  wire  _GEN_2199 = io_wb_info_i_4_valid & _GEN_2119 & _T_21 ? _GEN_2151 : _GEN_2095; // @[Rob.scala 283:75]
  wire  _GEN_2200 = io_wb_info_i_4_valid & _GEN_2119 & _T_21 ? _GEN_2152 : _GEN_2096; // @[Rob.scala 283:75]
  wire  _GEN_2201 = io_wb_info_i_4_valid & _GEN_2119 & _T_21 ? _GEN_2153 : _GEN_2097; // @[Rob.scala 283:75]
  wire  _GEN_2202 = io_wb_info_i_4_valid & _GEN_2119 & _T_21 ? _GEN_2154 : _GEN_2098; // @[Rob.scala 283:75]
  wire  _GEN_2203 = io_wb_info_i_4_valid & _GEN_2119 & _T_21 ? _GEN_2155 : _GEN_2099; // @[Rob.scala 283:75]
  wire  _GEN_2204 = io_wb_info_i_4_valid & _GEN_2119 & _T_21 ? _GEN_2156 : _GEN_2100; // @[Rob.scala 283:75]
  wire  _GEN_2205 = io_wb_info_i_4_valid & _GEN_2119 & _T_21 ? _GEN_2157 : _GEN_2101; // @[Rob.scala 283:75]
  wire  _GEN_2206 = io_wb_info_i_4_valid & _GEN_2119 & _T_21 ? _GEN_2158 : _GEN_2102; // @[Rob.scala 283:75]
  wire  _GEN_2207 = io_wb_info_i_4_valid & _GEN_2119 & _T_21 ? _GEN_2159 : _GEN_2103; // @[Rob.scala 283:75]
  wire [31:0] _GEN_2208 = io_wb_info_i_4_valid & _GEN_2119 & _T_21 ? _GEN_2160 : _GEN_2104; // @[Rob.scala 283:75]
  wire [31:0] _GEN_2209 = io_wb_info_i_4_valid & _GEN_2119 & _T_21 ? _GEN_2161 : _GEN_2105; // @[Rob.scala 283:75]
  wire [31:0] _GEN_2210 = io_wb_info_i_4_valid & _GEN_2119 & _T_21 ? _GEN_2162 : _GEN_2106; // @[Rob.scala 283:75]
  wire [31:0] _GEN_2211 = io_wb_info_i_4_valid & _GEN_2119 & _T_21 ? _GEN_2163 : _GEN_2107; // @[Rob.scala 283:75]
  wire [31:0] _GEN_2212 = io_wb_info_i_4_valid & _GEN_2119 & _T_21 ? _GEN_2164 : _GEN_2108; // @[Rob.scala 283:75]
  wire [31:0] _GEN_2213 = io_wb_info_i_4_valid & _GEN_2119 & _T_21 ? _GEN_2165 : _GEN_2109; // @[Rob.scala 283:75]
  wire [31:0] _GEN_2214 = io_wb_info_i_4_valid & _GEN_2119 & _T_21 ? _GEN_2166 : _GEN_2110; // @[Rob.scala 283:75]
  wire [31:0] _GEN_2215 = io_wb_info_i_4_valid & _GEN_2119 & _T_21 ? _GEN_2167 : _GEN_2111; // @[Rob.scala 283:75]
  wire  _init_op1_data_T = ~io_rob_init_info_bits_0_op1_in_rob; // @[Rob.scala 310:32]
  wire [31:0] _GEN_2217 = 3'h1 == io_rob_init_info_bits_0_op1_rob ? rob_info_1_commit_data : rob_info_0_commit_data; // @[Rob.scala 310:156 Rob.scala 310:156]
  wire [31:0] _GEN_2218 = 3'h2 == io_rob_init_info_bits_0_op1_rob ? rob_info_2_commit_data : _GEN_2217; // @[Rob.scala 310:156 Rob.scala 310:156]
  wire [31:0] _GEN_2219 = 3'h3 == io_rob_init_info_bits_0_op1_rob ? rob_info_3_commit_data : _GEN_2218; // @[Rob.scala 310:156 Rob.scala 310:156]
  wire [31:0] _GEN_2220 = 3'h4 == io_rob_init_info_bits_0_op1_rob ? rob_info_4_commit_data : _GEN_2219; // @[Rob.scala 310:156 Rob.scala 310:156]
  wire [31:0] _GEN_2221 = 3'h5 == io_rob_init_info_bits_0_op1_rob ? rob_info_5_commit_data : _GEN_2220; // @[Rob.scala 310:156 Rob.scala 310:156]
  wire [31:0] _GEN_2222 = 3'h6 == io_rob_init_info_bits_0_op1_rob ? rob_info_6_commit_data : _GEN_2221; // @[Rob.scala 310:156 Rob.scala 310:156]
  wire [31:0] _GEN_2223 = 3'h7 == io_rob_init_info_bits_0_op1_rob ? rob_info_7_commit_data : _GEN_2222; // @[Rob.scala 310:156 Rob.scala 310:156]
  reg [2:0] rob_commit_1_des_rob; // @[Rob.scala 341:23]
  reg  rob_commit_valid_1; // @[Rob.scala 342:33]
  reg [2:0] rob_commit_0_des_rob; // @[Rob.scala 341:23]
  reg  rob_commit_valid_0; // @[Rob.scala 342:33]
  wire  init_op1_hit_commit_0 = rob_commit_1_des_rob == io_rob_init_info_bits_0_op1_rob & rob_commit_valid_1 |
    rob_commit_0_des_rob == io_rob_init_info_bits_0_op1_rob & rob_commit_valid_0; // @[Rob.scala 359:92 Rob.scala 360:31]
  reg [31:0] rob_commit_1_commit_data; // @[Rob.scala 341:23]
  reg [31:0] rob_commit_0_commit_data; // @[Rob.scala 341:23]
  wire [31:0] _GEN_3473 = rob_commit_0_des_rob == io_rob_init_info_bits_0_op1_rob & rob_commit_valid_0 ?
    rob_commit_0_commit_data : 32'h0; // @[Rob.scala 359:92 Rob.scala 361:32]
  wire [31:0] init_op1_commit_data_0 = rob_commit_1_des_rob == io_rob_init_info_bits_0_op1_rob & rob_commit_valid_1 ?
    rob_commit_1_commit_data : _GEN_3473; // @[Rob.scala 359:92 Rob.scala 361:32]
  wire [31:0] _init_op1_data_T_1 = init_op1_hit_commit_0 ? init_op1_commit_data_0 : _GEN_2223; // @[Rob.scala 310:156]
  wire  init_op1_hit_wb_0 = io_wb_info_i_4_bits_rob_idx == io_rob_init_info_bits_0_op1_rob & io_wb_info_i_4_valid | (
    io_wb_info_i_3_bits_rob_idx == io_rob_init_info_bits_0_op1_rob & io_wb_info_i_3_valid | (io_wb_info_i_2_bits_rob_idx
     == io_rob_init_info_bits_0_op1_rob & io_wb_info_i_2_valid | (io_wb_info_i_1_bits_rob_idx ==
    io_rob_init_info_bits_0_op1_rob & io_wb_info_i_1_valid | io_wb_info_i_0_bits_rob_idx ==
    io_rob_init_info_bits_0_op1_rob & io_wb_info_i_0_valid))); // @[Rob.scala 371:101 Rob.scala 372:27]
  wire [31:0] _GEN_3489 = io_wb_info_i_0_bits_rob_idx == io_rob_init_info_bits_0_op1_rob & io_wb_info_i_0_valid ?
    io_wb_info_i_0_bits_data : 32'h0; // @[Rob.scala 371:101 Rob.scala 373:28]
  wire [31:0] _GEN_3493 = io_wb_info_i_1_bits_rob_idx == io_rob_init_info_bits_0_op1_rob & io_wb_info_i_1_valid ?
    io_wb_info_i_1_bits_data : _GEN_3489; // @[Rob.scala 371:101 Rob.scala 373:28]
  wire [31:0] _GEN_3497 = io_wb_info_i_2_bits_rob_idx == io_rob_init_info_bits_0_op1_rob & io_wb_info_i_2_valid ?
    io_wb_info_i_2_bits_data : _GEN_3493; // @[Rob.scala 371:101 Rob.scala 373:28]
  wire [31:0] _GEN_3501 = io_wb_info_i_3_bits_rob_idx == io_rob_init_info_bits_0_op1_rob & io_wb_info_i_3_valid ?
    io_wb_info_i_3_bits_data : _GEN_3497; // @[Rob.scala 371:101 Rob.scala 373:28]
  wire [31:0] init_op1_wb_data_0 = io_wb_info_i_4_bits_rob_idx == io_rob_init_info_bits_0_op1_rob & io_wb_info_i_4_valid
     ? io_wb_info_i_4_bits_data : _GEN_3501; // @[Rob.scala 371:101 Rob.scala 373:28]
  wire [31:0] _init_op1_data_T_2 = init_op1_hit_wb_0 ? init_op1_wb_data_0 : _init_op1_data_T_1; // @[Rob.scala 310:111]
  wire [31:0] init_op1_data = ~io_rob_init_info_bits_0_op1_in_rob ? io_rob_init_info_bits_0_op1_regData :
    _init_op1_data_T_2; // @[Rob.scala 310:31]
  wire  _init_op2_data_T = ~io_rob_init_info_bits_0_op2_in_rob; // @[Rob.scala 311:32]
  wire [31:0] _GEN_2225 = 3'h1 == io_rob_init_info_bits_0_op2_rob ? rob_info_1_commit_data : rob_info_0_commit_data; // @[Rob.scala 311:156 Rob.scala 311:156]
  wire [31:0] _GEN_2226 = 3'h2 == io_rob_init_info_bits_0_op2_rob ? rob_info_2_commit_data : _GEN_2225; // @[Rob.scala 311:156 Rob.scala 311:156]
  wire [31:0] _GEN_2227 = 3'h3 == io_rob_init_info_bits_0_op2_rob ? rob_info_3_commit_data : _GEN_2226; // @[Rob.scala 311:156 Rob.scala 311:156]
  wire [31:0] _GEN_2228 = 3'h4 == io_rob_init_info_bits_0_op2_rob ? rob_info_4_commit_data : _GEN_2227; // @[Rob.scala 311:156 Rob.scala 311:156]
  wire [31:0] _GEN_2229 = 3'h5 == io_rob_init_info_bits_0_op2_rob ? rob_info_5_commit_data : _GEN_2228; // @[Rob.scala 311:156 Rob.scala 311:156]
  wire [31:0] _GEN_2230 = 3'h6 == io_rob_init_info_bits_0_op2_rob ? rob_info_6_commit_data : _GEN_2229; // @[Rob.scala 311:156 Rob.scala 311:156]
  wire [31:0] _GEN_2231 = 3'h7 == io_rob_init_info_bits_0_op2_rob ? rob_info_7_commit_data : _GEN_2230; // @[Rob.scala 311:156 Rob.scala 311:156]
  wire  init_op2_hit_commit_0 = rob_commit_1_des_rob == io_rob_init_info_bits_0_op2_rob & rob_commit_valid_1 |
    rob_commit_0_des_rob == io_rob_init_info_bits_0_op2_rob & rob_commit_valid_0; // @[Rob.scala 363:92 Rob.scala 364:31]
  wire [31:0] _GEN_3475 = rob_commit_0_des_rob == io_rob_init_info_bits_0_op2_rob & rob_commit_valid_0 ?
    rob_commit_0_commit_data : 32'h0; // @[Rob.scala 363:92 Rob.scala 365:32]
  wire [31:0] init_op2_commit_data_0 = rob_commit_1_des_rob == io_rob_init_info_bits_0_op2_rob & rob_commit_valid_1 ?
    rob_commit_1_commit_data : _GEN_3475; // @[Rob.scala 363:92 Rob.scala 365:32]
  wire [31:0] _init_op2_data_T_1 = init_op2_hit_commit_0 ? init_op2_commit_data_0 : _GEN_2231; // @[Rob.scala 311:156]
  wire  init_op2_hit_wb_0 = io_wb_info_i_4_bits_rob_idx == io_rob_init_info_bits_0_op2_rob & io_wb_info_i_4_valid | (
    io_wb_info_i_3_bits_rob_idx == io_rob_init_info_bits_0_op2_rob & io_wb_info_i_3_valid | (io_wb_info_i_2_bits_rob_idx
     == io_rob_init_info_bits_0_op2_rob & io_wb_info_i_2_valid | (io_wb_info_i_1_bits_rob_idx ==
    io_rob_init_info_bits_0_op2_rob & io_wb_info_i_1_valid | io_wb_info_i_0_bits_rob_idx ==
    io_rob_init_info_bits_0_op2_rob & io_wb_info_i_0_valid))); // @[Rob.scala 375:101 Rob.scala 376:27]
  wire [31:0] _GEN_3491 = io_wb_info_i_0_bits_rob_idx == io_rob_init_info_bits_0_op2_rob & io_wb_info_i_0_valid ?
    io_wb_info_i_0_bits_data : 32'h0; // @[Rob.scala 375:101 Rob.scala 377:28]
  wire [31:0] _GEN_3495 = io_wb_info_i_1_bits_rob_idx == io_rob_init_info_bits_0_op2_rob & io_wb_info_i_1_valid ?
    io_wb_info_i_1_bits_data : _GEN_3491; // @[Rob.scala 375:101 Rob.scala 377:28]
  wire [31:0] _GEN_3499 = io_wb_info_i_2_bits_rob_idx == io_rob_init_info_bits_0_op2_rob & io_wb_info_i_2_valid ?
    io_wb_info_i_2_bits_data : _GEN_3495; // @[Rob.scala 375:101 Rob.scala 377:28]
  wire [31:0] _GEN_3503 = io_wb_info_i_3_bits_rob_idx == io_rob_init_info_bits_0_op2_rob & io_wb_info_i_3_valid ?
    io_wb_info_i_3_bits_data : _GEN_3499; // @[Rob.scala 375:101 Rob.scala 377:28]
  wire [31:0] init_op2_wb_data_0 = io_wb_info_i_4_bits_rob_idx == io_rob_init_info_bits_0_op2_rob & io_wb_info_i_4_valid
     ? io_wb_info_i_4_bits_data : _GEN_3503; // @[Rob.scala 375:101 Rob.scala 377:28]
  wire [31:0] _init_op2_data_T_2 = init_op2_hit_wb_0 ? init_op2_wb_data_0 : _init_op2_data_T_1; // @[Rob.scala 311:111]
  wire [31:0] init_op2_data = ~io_rob_init_info_bits_0_op2_in_rob ? io_rob_init_info_bits_0_op2_regData :
    _init_op2_data_T_2; // @[Rob.scala 311:31]
  wire  _GEN_2233 = 3'h1 == io_rob_init_info_bits_0_op1_rob ? rob_info_1_commit_ready : rob_info_0_commit_ready; // @[Rob.scala 312:59 Rob.scala 312:59]
  wire  _GEN_2234 = 3'h2 == io_rob_init_info_bits_0_op1_rob ? rob_info_2_commit_ready : _GEN_2233; // @[Rob.scala 312:59 Rob.scala 312:59]
  wire  _GEN_2235 = 3'h3 == io_rob_init_info_bits_0_op1_rob ? rob_info_3_commit_ready : _GEN_2234; // @[Rob.scala 312:59 Rob.scala 312:59]
  wire  _GEN_2236 = 3'h4 == io_rob_init_info_bits_0_op1_rob ? rob_info_4_commit_ready : _GEN_2235; // @[Rob.scala 312:59 Rob.scala 312:59]
  wire  _GEN_2237 = 3'h5 == io_rob_init_info_bits_0_op1_rob ? rob_info_5_commit_ready : _GEN_2236; // @[Rob.scala 312:59 Rob.scala 312:59]
  wire  _GEN_2238 = 3'h6 == io_rob_init_info_bits_0_op1_rob ? rob_info_6_commit_ready : _GEN_2237; // @[Rob.scala 312:59 Rob.scala 312:59]
  wire  _GEN_2239 = 3'h7 == io_rob_init_info_bits_0_op1_rob ? rob_info_7_commit_ready : _GEN_2238; // @[Rob.scala 312:59 Rob.scala 312:59]
  wire  _GEN_2241 = 3'h1 == io_rob_init_info_bits_0_op1_rob ? rob_info_1_is_valid : rob_info_0_is_valid; // @[Rob.scala 312:59 Rob.scala 312:59]
  wire  _GEN_2242 = 3'h2 == io_rob_init_info_bits_0_op1_rob ? rob_info_2_is_valid : _GEN_2241; // @[Rob.scala 312:59 Rob.scala 312:59]
  wire  _GEN_2243 = 3'h3 == io_rob_init_info_bits_0_op1_rob ? rob_info_3_is_valid : _GEN_2242; // @[Rob.scala 312:59 Rob.scala 312:59]
  wire  _GEN_2244 = 3'h4 == io_rob_init_info_bits_0_op1_rob ? rob_info_4_is_valid : _GEN_2243; // @[Rob.scala 312:59 Rob.scala 312:59]
  wire  _GEN_2245 = 3'h5 == io_rob_init_info_bits_0_op1_rob ? rob_info_5_is_valid : _GEN_2244; // @[Rob.scala 312:59 Rob.scala 312:59]
  wire  _GEN_2246 = 3'h6 == io_rob_init_info_bits_0_op1_rob ? rob_info_6_is_valid : _GEN_2245; // @[Rob.scala 312:59 Rob.scala 312:59]
  wire  _GEN_2247 = 3'h7 == io_rob_init_info_bits_0_op1_rob ? rob_info_7_is_valid : _GEN_2246; // @[Rob.scala 312:59 Rob.scala 312:59]
  wire  init_op1_hit_rob = _GEN_2239 & _GEN_2247 | init_op1_hit_wb_0 | init_op1_hit_commit_0; // @[Rob.scala 312:111]
  wire  _GEN_2249 = 3'h1 == io_rob_init_info_bits_0_op2_rob ? rob_info_1_commit_ready : rob_info_0_commit_ready; // @[Rob.scala 313:59 Rob.scala 313:59]
  wire  _GEN_2250 = 3'h2 == io_rob_init_info_bits_0_op2_rob ? rob_info_2_commit_ready : _GEN_2249; // @[Rob.scala 313:59 Rob.scala 313:59]
  wire  _GEN_2251 = 3'h3 == io_rob_init_info_bits_0_op2_rob ? rob_info_3_commit_ready : _GEN_2250; // @[Rob.scala 313:59 Rob.scala 313:59]
  wire  _GEN_2252 = 3'h4 == io_rob_init_info_bits_0_op2_rob ? rob_info_4_commit_ready : _GEN_2251; // @[Rob.scala 313:59 Rob.scala 313:59]
  wire  _GEN_2253 = 3'h5 == io_rob_init_info_bits_0_op2_rob ? rob_info_5_commit_ready : _GEN_2252; // @[Rob.scala 313:59 Rob.scala 313:59]
  wire  _GEN_2254 = 3'h6 == io_rob_init_info_bits_0_op2_rob ? rob_info_6_commit_ready : _GEN_2253; // @[Rob.scala 313:59 Rob.scala 313:59]
  wire  _GEN_2255 = 3'h7 == io_rob_init_info_bits_0_op2_rob ? rob_info_7_commit_ready : _GEN_2254; // @[Rob.scala 313:59 Rob.scala 313:59]
  wire  _GEN_2257 = 3'h1 == io_rob_init_info_bits_0_op2_rob ? rob_info_1_is_valid : rob_info_0_is_valid; // @[Rob.scala 313:59 Rob.scala 313:59]
  wire  _GEN_2258 = 3'h2 == io_rob_init_info_bits_0_op2_rob ? rob_info_2_is_valid : _GEN_2257; // @[Rob.scala 313:59 Rob.scala 313:59]
  wire  _GEN_2259 = 3'h3 == io_rob_init_info_bits_0_op2_rob ? rob_info_3_is_valid : _GEN_2258; // @[Rob.scala 313:59 Rob.scala 313:59]
  wire  _GEN_2260 = 3'h4 == io_rob_init_info_bits_0_op2_rob ? rob_info_4_is_valid : _GEN_2259; // @[Rob.scala 313:59 Rob.scala 313:59]
  wire  _GEN_2261 = 3'h5 == io_rob_init_info_bits_0_op2_rob ? rob_info_5_is_valid : _GEN_2260; // @[Rob.scala 313:59 Rob.scala 313:59]
  wire  _GEN_2262 = 3'h6 == io_rob_init_info_bits_0_op2_rob ? rob_info_6_is_valid : _GEN_2261; // @[Rob.scala 313:59 Rob.scala 313:59]
  wire  _GEN_2263 = 3'h7 == io_rob_init_info_bits_0_op2_rob ? rob_info_7_is_valid : _GEN_2262; // @[Rob.scala 313:59 Rob.scala 313:59]
  wire  init_op2_hit_rob = _GEN_2255 & _GEN_2263 | init_op2_hit_wb_0 | init_op2_hit_commit_0; // @[Rob.scala 313:111]
  wire [31:0] _GEN_2264 = 3'h0 == io_rob_init_info_bits_0_des_rob ? init_op1_data : _GEN_1552; // @[Rob.scala 316:34 Rob.scala 316:34]
  wire [31:0] _GEN_2265 = 3'h1 == io_rob_init_info_bits_0_des_rob ? init_op1_data : _GEN_1572; // @[Rob.scala 316:34 Rob.scala 316:34]
  wire [31:0] _GEN_2266 = 3'h2 == io_rob_init_info_bits_0_des_rob ? init_op1_data : _GEN_1592; // @[Rob.scala 316:34 Rob.scala 316:34]
  wire [31:0] _GEN_2267 = 3'h3 == io_rob_init_info_bits_0_des_rob ? init_op1_data : _GEN_1612; // @[Rob.scala 316:34 Rob.scala 316:34]
  wire [31:0] _GEN_2268 = 3'h4 == io_rob_init_info_bits_0_des_rob ? init_op1_data : _GEN_1632; // @[Rob.scala 316:34 Rob.scala 316:34]
  wire [31:0] _GEN_2269 = 3'h5 == io_rob_init_info_bits_0_des_rob ? init_op1_data : _GEN_1652; // @[Rob.scala 316:34 Rob.scala 316:34]
  wire [31:0] _GEN_2270 = 3'h6 == io_rob_init_info_bits_0_des_rob ? init_op1_data : _GEN_1672; // @[Rob.scala 316:34 Rob.scala 316:34]
  wire [31:0] _GEN_2271 = 3'h7 == io_rob_init_info_bits_0_des_rob ? init_op1_data : _GEN_1692; // @[Rob.scala 316:34 Rob.scala 316:34]
  wire [31:0] _GEN_2272 = 3'h0 == io_rob_init_info_bits_0_des_rob ? init_op2_data : _GEN_1554; // @[Rob.scala 317:34 Rob.scala 317:34]
  wire [31:0] _GEN_2273 = 3'h1 == io_rob_init_info_bits_0_des_rob ? init_op2_data : _GEN_1574; // @[Rob.scala 317:34 Rob.scala 317:34]
  wire [31:0] _GEN_2274 = 3'h2 == io_rob_init_info_bits_0_des_rob ? init_op2_data : _GEN_1594; // @[Rob.scala 317:34 Rob.scala 317:34]
  wire [31:0] _GEN_2275 = 3'h3 == io_rob_init_info_bits_0_des_rob ? init_op2_data : _GEN_1614; // @[Rob.scala 317:34 Rob.scala 317:34]
  wire [31:0] _GEN_2276 = 3'h4 == io_rob_init_info_bits_0_des_rob ? init_op2_data : _GEN_1634; // @[Rob.scala 317:34 Rob.scala 317:34]
  wire [31:0] _GEN_2277 = 3'h5 == io_rob_init_info_bits_0_des_rob ? init_op2_data : _GEN_1654; // @[Rob.scala 317:34 Rob.scala 317:34]
  wire [31:0] _GEN_2278 = 3'h6 == io_rob_init_info_bits_0_des_rob ? init_op2_data : _GEN_1674; // @[Rob.scala 317:34 Rob.scala 317:34]
  wire [31:0] _GEN_2279 = 3'h7 == io_rob_init_info_bits_0_des_rob ? init_op2_data : _GEN_1694; // @[Rob.scala 317:34 Rob.scala 317:34]
  wire [2:0] _GEN_2280 = 3'h0 == io_rob_init_info_bits_0_des_rob ? io_rob_init_info_bits_0_op1_rob : rob_info_0_op1_tag; // @[Rob.scala 318:33 Rob.scala 318:33 Rob.scala 175:27]
  wire [2:0] _GEN_2281 = 3'h1 == io_rob_init_info_bits_0_des_rob ? io_rob_init_info_bits_0_op1_rob : rob_info_1_op1_tag; // @[Rob.scala 318:33 Rob.scala 318:33 Rob.scala 175:27]
  wire [2:0] _GEN_2282 = 3'h2 == io_rob_init_info_bits_0_des_rob ? io_rob_init_info_bits_0_op1_rob : rob_info_2_op1_tag; // @[Rob.scala 318:33 Rob.scala 318:33 Rob.scala 175:27]
  wire [2:0] _GEN_2283 = 3'h3 == io_rob_init_info_bits_0_des_rob ? io_rob_init_info_bits_0_op1_rob : rob_info_3_op1_tag; // @[Rob.scala 318:33 Rob.scala 318:33 Rob.scala 175:27]
  wire [2:0] _GEN_2284 = 3'h4 == io_rob_init_info_bits_0_des_rob ? io_rob_init_info_bits_0_op1_rob : rob_info_4_op1_tag; // @[Rob.scala 318:33 Rob.scala 318:33 Rob.scala 175:27]
  wire [2:0] _GEN_2285 = 3'h5 == io_rob_init_info_bits_0_des_rob ? io_rob_init_info_bits_0_op1_rob : rob_info_5_op1_tag; // @[Rob.scala 318:33 Rob.scala 318:33 Rob.scala 175:27]
  wire [2:0] _GEN_2286 = 3'h6 == io_rob_init_info_bits_0_des_rob ? io_rob_init_info_bits_0_op1_rob : rob_info_6_op1_tag; // @[Rob.scala 318:33 Rob.scala 318:33 Rob.scala 175:27]
  wire [2:0] _GEN_2287 = 3'h7 == io_rob_init_info_bits_0_des_rob ? io_rob_init_info_bits_0_op1_rob : rob_info_7_op1_tag; // @[Rob.scala 318:33 Rob.scala 318:33 Rob.scala 175:27]
  wire [2:0] _GEN_2288 = 3'h0 == io_rob_init_info_bits_0_des_rob ? io_rob_init_info_bits_0_op2_rob : rob_info_0_op2_tag; // @[Rob.scala 319:33 Rob.scala 319:33 Rob.scala 175:27]
  wire [2:0] _GEN_2289 = 3'h1 == io_rob_init_info_bits_0_des_rob ? io_rob_init_info_bits_0_op2_rob : rob_info_1_op2_tag; // @[Rob.scala 319:33 Rob.scala 319:33 Rob.scala 175:27]
  wire [2:0] _GEN_2290 = 3'h2 == io_rob_init_info_bits_0_des_rob ? io_rob_init_info_bits_0_op2_rob : rob_info_2_op2_tag; // @[Rob.scala 319:33 Rob.scala 319:33 Rob.scala 175:27]
  wire [2:0] _GEN_2291 = 3'h3 == io_rob_init_info_bits_0_des_rob ? io_rob_init_info_bits_0_op2_rob : rob_info_3_op2_tag; // @[Rob.scala 319:33 Rob.scala 319:33 Rob.scala 175:27]
  wire [2:0] _GEN_2292 = 3'h4 == io_rob_init_info_bits_0_des_rob ? io_rob_init_info_bits_0_op2_rob : rob_info_4_op2_tag; // @[Rob.scala 319:33 Rob.scala 319:33 Rob.scala 175:27]
  wire [2:0] _GEN_2293 = 3'h5 == io_rob_init_info_bits_0_des_rob ? io_rob_init_info_bits_0_op2_rob : rob_info_5_op2_tag; // @[Rob.scala 319:33 Rob.scala 319:33 Rob.scala 175:27]
  wire [2:0] _GEN_2294 = 3'h6 == io_rob_init_info_bits_0_des_rob ? io_rob_init_info_bits_0_op2_rob : rob_info_6_op2_tag; // @[Rob.scala 319:33 Rob.scala 319:33 Rob.scala 175:27]
  wire [2:0] _GEN_2295 = 3'h7 == io_rob_init_info_bits_0_des_rob ? io_rob_init_info_bits_0_op2_rob : rob_info_7_op2_tag; // @[Rob.scala 319:33 Rob.scala 319:33 Rob.scala 175:27]
  wire  _GEN_2296 = 3'h0 == io_rob_init_info_bits_0_des_rob ? _init_op1_data_T | init_op1_hit_rob : _GEN_1553; // @[Rob.scala 320:35 Rob.scala 320:35]
  wire  _GEN_2297 = 3'h1 == io_rob_init_info_bits_0_des_rob ? _init_op1_data_T | init_op1_hit_rob : _GEN_1573; // @[Rob.scala 320:35 Rob.scala 320:35]
  wire  _GEN_2298 = 3'h2 == io_rob_init_info_bits_0_des_rob ? _init_op1_data_T | init_op1_hit_rob : _GEN_1593; // @[Rob.scala 320:35 Rob.scala 320:35]
  wire  _GEN_2299 = 3'h3 == io_rob_init_info_bits_0_des_rob ? _init_op1_data_T | init_op1_hit_rob : _GEN_1613; // @[Rob.scala 320:35 Rob.scala 320:35]
  wire  _GEN_2300 = 3'h4 == io_rob_init_info_bits_0_des_rob ? _init_op1_data_T | init_op1_hit_rob : _GEN_1633; // @[Rob.scala 320:35 Rob.scala 320:35]
  wire  _GEN_2301 = 3'h5 == io_rob_init_info_bits_0_des_rob ? _init_op1_data_T | init_op1_hit_rob : _GEN_1653; // @[Rob.scala 320:35 Rob.scala 320:35]
  wire  _GEN_2302 = 3'h6 == io_rob_init_info_bits_0_des_rob ? _init_op1_data_T | init_op1_hit_rob : _GEN_1673; // @[Rob.scala 320:35 Rob.scala 320:35]
  wire  _GEN_2303 = 3'h7 == io_rob_init_info_bits_0_des_rob ? _init_op1_data_T | init_op1_hit_rob : _GEN_1693; // @[Rob.scala 320:35 Rob.scala 320:35]
  wire  _GEN_2304 = 3'h0 == io_rob_init_info_bits_0_des_rob ? _init_op2_data_T | init_op2_hit_rob : _GEN_1555; // @[Rob.scala 321:35 Rob.scala 321:35]
  wire  _GEN_2305 = 3'h1 == io_rob_init_info_bits_0_des_rob ? _init_op2_data_T | init_op2_hit_rob : _GEN_1575; // @[Rob.scala 321:35 Rob.scala 321:35]
  wire  _GEN_2306 = 3'h2 == io_rob_init_info_bits_0_des_rob ? _init_op2_data_T | init_op2_hit_rob : _GEN_1595; // @[Rob.scala 321:35 Rob.scala 321:35]
  wire  _GEN_2307 = 3'h3 == io_rob_init_info_bits_0_des_rob ? _init_op2_data_T | init_op2_hit_rob : _GEN_1615; // @[Rob.scala 321:35 Rob.scala 321:35]
  wire  _GEN_2308 = 3'h4 == io_rob_init_info_bits_0_des_rob ? _init_op2_data_T | init_op2_hit_rob : _GEN_1635; // @[Rob.scala 321:35 Rob.scala 321:35]
  wire  _GEN_2309 = 3'h5 == io_rob_init_info_bits_0_des_rob ? _init_op2_data_T | init_op2_hit_rob : _GEN_1655; // @[Rob.scala 321:35 Rob.scala 321:35]
  wire  _GEN_2310 = 3'h6 == io_rob_init_info_bits_0_des_rob ? _init_op2_data_T | init_op2_hit_rob : _GEN_1675; // @[Rob.scala 321:35 Rob.scala 321:35]
  wire  _GEN_2311 = 3'h7 == io_rob_init_info_bits_0_des_rob ? _init_op2_data_T | init_op2_hit_rob : _GEN_1695; // @[Rob.scala 321:35 Rob.scala 321:35]
  wire  _GEN_2312 = 3'h0 == io_rob_init_info_bits_0_des_rob | _GEN_1424; // @[Rob.scala 322:33 Rob.scala 322:33]
  wire  _GEN_2313 = 3'h1 == io_rob_init_info_bits_0_des_rob | _GEN_1425; // @[Rob.scala 322:33 Rob.scala 322:33]
  wire  _GEN_2314 = 3'h2 == io_rob_init_info_bits_0_des_rob | _GEN_1426; // @[Rob.scala 322:33 Rob.scala 322:33]
  wire  _GEN_2315 = 3'h3 == io_rob_init_info_bits_0_des_rob | _GEN_1427; // @[Rob.scala 322:33 Rob.scala 322:33]
  wire  _GEN_2316 = 3'h4 == io_rob_init_info_bits_0_des_rob | _GEN_1428; // @[Rob.scala 322:33 Rob.scala 322:33]
  wire  _GEN_2317 = 3'h5 == io_rob_init_info_bits_0_des_rob | _GEN_1429; // @[Rob.scala 322:33 Rob.scala 322:33]
  wire  _GEN_2318 = 3'h6 == io_rob_init_info_bits_0_des_rob | _GEN_1430; // @[Rob.scala 322:33 Rob.scala 322:33]
  wire  _GEN_2319 = 3'h7 == io_rob_init_info_bits_0_des_rob | _GEN_1431; // @[Rob.scala 322:33 Rob.scala 322:33]
  wire [31:0] _GEN_2320 = io_rob_init_info_valid & io_rob_init_info_bits_0_is_valid & _T_21 ? _GEN_2264 : _GEN_1552; // @[Rob.scala 315:86]
  wire [31:0] _GEN_2321 = io_rob_init_info_valid & io_rob_init_info_bits_0_is_valid & _T_21 ? _GEN_2265 : _GEN_1572; // @[Rob.scala 315:86]
  wire [31:0] _GEN_2322 = io_rob_init_info_valid & io_rob_init_info_bits_0_is_valid & _T_21 ? _GEN_2266 : _GEN_1592; // @[Rob.scala 315:86]
  wire [31:0] _GEN_2323 = io_rob_init_info_valid & io_rob_init_info_bits_0_is_valid & _T_21 ? _GEN_2267 : _GEN_1612; // @[Rob.scala 315:86]
  wire [31:0] _GEN_2324 = io_rob_init_info_valid & io_rob_init_info_bits_0_is_valid & _T_21 ? _GEN_2268 : _GEN_1632; // @[Rob.scala 315:86]
  wire [31:0] _GEN_2325 = io_rob_init_info_valid & io_rob_init_info_bits_0_is_valid & _T_21 ? _GEN_2269 : _GEN_1652; // @[Rob.scala 315:86]
  wire [31:0] _GEN_2326 = io_rob_init_info_valid & io_rob_init_info_bits_0_is_valid & _T_21 ? _GEN_2270 : _GEN_1672; // @[Rob.scala 315:86]
  wire [31:0] _GEN_2327 = io_rob_init_info_valid & io_rob_init_info_bits_0_is_valid & _T_21 ? _GEN_2271 : _GEN_1692; // @[Rob.scala 315:86]
  wire [31:0] _GEN_2328 = io_rob_init_info_valid & io_rob_init_info_bits_0_is_valid & _T_21 ? _GEN_2272 : _GEN_1554; // @[Rob.scala 315:86]
  wire [31:0] _GEN_2329 = io_rob_init_info_valid & io_rob_init_info_bits_0_is_valid & _T_21 ? _GEN_2273 : _GEN_1574; // @[Rob.scala 315:86]
  wire [31:0] _GEN_2330 = io_rob_init_info_valid & io_rob_init_info_bits_0_is_valid & _T_21 ? _GEN_2274 : _GEN_1594; // @[Rob.scala 315:86]
  wire [31:0] _GEN_2331 = io_rob_init_info_valid & io_rob_init_info_bits_0_is_valid & _T_21 ? _GEN_2275 : _GEN_1614; // @[Rob.scala 315:86]
  wire [31:0] _GEN_2332 = io_rob_init_info_valid & io_rob_init_info_bits_0_is_valid & _T_21 ? _GEN_2276 : _GEN_1634; // @[Rob.scala 315:86]
  wire [31:0] _GEN_2333 = io_rob_init_info_valid & io_rob_init_info_bits_0_is_valid & _T_21 ? _GEN_2277 : _GEN_1654; // @[Rob.scala 315:86]
  wire [31:0] _GEN_2334 = io_rob_init_info_valid & io_rob_init_info_bits_0_is_valid & _T_21 ? _GEN_2278 : _GEN_1674; // @[Rob.scala 315:86]
  wire [31:0] _GEN_2335 = io_rob_init_info_valid & io_rob_init_info_bits_0_is_valid & _T_21 ? _GEN_2279 : _GEN_1694; // @[Rob.scala 315:86]
  wire [2:0] _GEN_2336 = io_rob_init_info_valid & io_rob_init_info_bits_0_is_valid & _T_21 ? _GEN_2280 :
    rob_info_0_op1_tag; // @[Rob.scala 315:86 Rob.scala 175:27]
  wire [2:0] _GEN_2337 = io_rob_init_info_valid & io_rob_init_info_bits_0_is_valid & _T_21 ? _GEN_2281 :
    rob_info_1_op1_tag; // @[Rob.scala 315:86 Rob.scala 175:27]
  wire [2:0] _GEN_2338 = io_rob_init_info_valid & io_rob_init_info_bits_0_is_valid & _T_21 ? _GEN_2282 :
    rob_info_2_op1_tag; // @[Rob.scala 315:86 Rob.scala 175:27]
  wire [2:0] _GEN_2339 = io_rob_init_info_valid & io_rob_init_info_bits_0_is_valid & _T_21 ? _GEN_2283 :
    rob_info_3_op1_tag; // @[Rob.scala 315:86 Rob.scala 175:27]
  wire [2:0] _GEN_2340 = io_rob_init_info_valid & io_rob_init_info_bits_0_is_valid & _T_21 ? _GEN_2284 :
    rob_info_4_op1_tag; // @[Rob.scala 315:86 Rob.scala 175:27]
  wire [2:0] _GEN_2341 = io_rob_init_info_valid & io_rob_init_info_bits_0_is_valid & _T_21 ? _GEN_2285 :
    rob_info_5_op1_tag; // @[Rob.scala 315:86 Rob.scala 175:27]
  wire [2:0] _GEN_2342 = io_rob_init_info_valid & io_rob_init_info_bits_0_is_valid & _T_21 ? _GEN_2286 :
    rob_info_6_op1_tag; // @[Rob.scala 315:86 Rob.scala 175:27]
  wire [2:0] _GEN_2343 = io_rob_init_info_valid & io_rob_init_info_bits_0_is_valid & _T_21 ? _GEN_2287 :
    rob_info_7_op1_tag; // @[Rob.scala 315:86 Rob.scala 175:27]
  wire [2:0] _GEN_2344 = io_rob_init_info_valid & io_rob_init_info_bits_0_is_valid & _T_21 ? _GEN_2288 :
    rob_info_0_op2_tag; // @[Rob.scala 315:86 Rob.scala 175:27]
  wire [2:0] _GEN_2345 = io_rob_init_info_valid & io_rob_init_info_bits_0_is_valid & _T_21 ? _GEN_2289 :
    rob_info_1_op2_tag; // @[Rob.scala 315:86 Rob.scala 175:27]
  wire [2:0] _GEN_2346 = io_rob_init_info_valid & io_rob_init_info_bits_0_is_valid & _T_21 ? _GEN_2290 :
    rob_info_2_op2_tag; // @[Rob.scala 315:86 Rob.scala 175:27]
  wire [2:0] _GEN_2347 = io_rob_init_info_valid & io_rob_init_info_bits_0_is_valid & _T_21 ? _GEN_2291 :
    rob_info_3_op2_tag; // @[Rob.scala 315:86 Rob.scala 175:27]
  wire [2:0] _GEN_2348 = io_rob_init_info_valid & io_rob_init_info_bits_0_is_valid & _T_21 ? _GEN_2292 :
    rob_info_4_op2_tag; // @[Rob.scala 315:86 Rob.scala 175:27]
  wire [2:0] _GEN_2349 = io_rob_init_info_valid & io_rob_init_info_bits_0_is_valid & _T_21 ? _GEN_2293 :
    rob_info_5_op2_tag; // @[Rob.scala 315:86 Rob.scala 175:27]
  wire [2:0] _GEN_2350 = io_rob_init_info_valid & io_rob_init_info_bits_0_is_valid & _T_21 ? _GEN_2294 :
    rob_info_6_op2_tag; // @[Rob.scala 315:86 Rob.scala 175:27]
  wire [2:0] _GEN_2351 = io_rob_init_info_valid & io_rob_init_info_bits_0_is_valid & _T_21 ? _GEN_2295 :
    rob_info_7_op2_tag; // @[Rob.scala 315:86 Rob.scala 175:27]
  wire  _GEN_2352 = io_rob_init_info_valid & io_rob_init_info_bits_0_is_valid & _T_21 ? _GEN_2296 : _GEN_1553; // @[Rob.scala 315:86]
  wire  _GEN_2353 = io_rob_init_info_valid & io_rob_init_info_bits_0_is_valid & _T_21 ? _GEN_2297 : _GEN_1573; // @[Rob.scala 315:86]
  wire  _GEN_2354 = io_rob_init_info_valid & io_rob_init_info_bits_0_is_valid & _T_21 ? _GEN_2298 : _GEN_1593; // @[Rob.scala 315:86]
  wire  _GEN_2355 = io_rob_init_info_valid & io_rob_init_info_bits_0_is_valid & _T_21 ? _GEN_2299 : _GEN_1613; // @[Rob.scala 315:86]
  wire  _GEN_2356 = io_rob_init_info_valid & io_rob_init_info_bits_0_is_valid & _T_21 ? _GEN_2300 : _GEN_1633; // @[Rob.scala 315:86]
  wire  _GEN_2357 = io_rob_init_info_valid & io_rob_init_info_bits_0_is_valid & _T_21 ? _GEN_2301 : _GEN_1653; // @[Rob.scala 315:86]
  wire  _GEN_2358 = io_rob_init_info_valid & io_rob_init_info_bits_0_is_valid & _T_21 ? _GEN_2302 : _GEN_1673; // @[Rob.scala 315:86]
  wire  _GEN_2359 = io_rob_init_info_valid & io_rob_init_info_bits_0_is_valid & _T_21 ? _GEN_2303 : _GEN_1693; // @[Rob.scala 315:86]
  wire  _GEN_2360 = io_rob_init_info_valid & io_rob_init_info_bits_0_is_valid & _T_21 ? _GEN_2304 : _GEN_1555; // @[Rob.scala 315:86]
  wire  _GEN_2361 = io_rob_init_info_valid & io_rob_init_info_bits_0_is_valid & _T_21 ? _GEN_2305 : _GEN_1575; // @[Rob.scala 315:86]
  wire  _GEN_2362 = io_rob_init_info_valid & io_rob_init_info_bits_0_is_valid & _T_21 ? _GEN_2306 : _GEN_1595; // @[Rob.scala 315:86]
  wire  _GEN_2363 = io_rob_init_info_valid & io_rob_init_info_bits_0_is_valid & _T_21 ? _GEN_2307 : _GEN_1615; // @[Rob.scala 315:86]
  wire  _GEN_2364 = io_rob_init_info_valid & io_rob_init_info_bits_0_is_valid & _T_21 ? _GEN_2308 : _GEN_1635; // @[Rob.scala 315:86]
  wire  _GEN_2365 = io_rob_init_info_valid & io_rob_init_info_bits_0_is_valid & _T_21 ? _GEN_2309 : _GEN_1655; // @[Rob.scala 315:86]
  wire  _GEN_2366 = io_rob_init_info_valid & io_rob_init_info_bits_0_is_valid & _T_21 ? _GEN_2310 : _GEN_1675; // @[Rob.scala 315:86]
  wire  _GEN_2367 = io_rob_init_info_valid & io_rob_init_info_bits_0_is_valid & _T_21 ? _GEN_2311 : _GEN_1695; // @[Rob.scala 315:86]
  wire  _GEN_2368 = io_rob_init_info_valid & io_rob_init_info_bits_0_is_valid & _T_21 ? _GEN_2312 : _GEN_1424; // @[Rob.scala 315:86]
  wire  _GEN_2369 = io_rob_init_info_valid & io_rob_init_info_bits_0_is_valid & _T_21 ? _GEN_2313 : _GEN_1425; // @[Rob.scala 315:86]
  wire  _GEN_2370 = io_rob_init_info_valid & io_rob_init_info_bits_0_is_valid & _T_21 ? _GEN_2314 : _GEN_1426; // @[Rob.scala 315:86]
  wire  _GEN_2371 = io_rob_init_info_valid & io_rob_init_info_bits_0_is_valid & _T_21 ? _GEN_2315 : _GEN_1427; // @[Rob.scala 315:86]
  wire  _GEN_2372 = io_rob_init_info_valid & io_rob_init_info_bits_0_is_valid & _T_21 ? _GEN_2316 : _GEN_1428; // @[Rob.scala 315:86]
  wire  _GEN_2373 = io_rob_init_info_valid & io_rob_init_info_bits_0_is_valid & _T_21 ? _GEN_2317 : _GEN_1429; // @[Rob.scala 315:86]
  wire  _GEN_2374 = io_rob_init_info_valid & io_rob_init_info_bits_0_is_valid & _T_21 ? _GEN_2318 : _GEN_1430; // @[Rob.scala 315:86]
  wire  _GEN_2375 = io_rob_init_info_valid & io_rob_init_info_bits_0_is_valid & _T_21 ? _GEN_2319 : _GEN_1431; // @[Rob.scala 315:86]
  wire  _init_op1_data_T_3 = ~io_rob_init_info_bits_1_op1_in_rob; // @[Rob.scala 310:32]
  wire [31:0] _GEN_2377 = 3'h1 == io_rob_init_info_bits_1_op1_rob ? rob_info_1_commit_data : rob_info_0_commit_data; // @[Rob.scala 310:156 Rob.scala 310:156]
  wire [31:0] _GEN_2378 = 3'h2 == io_rob_init_info_bits_1_op1_rob ? rob_info_2_commit_data : _GEN_2377; // @[Rob.scala 310:156 Rob.scala 310:156]
  wire [31:0] _GEN_2379 = 3'h3 == io_rob_init_info_bits_1_op1_rob ? rob_info_3_commit_data : _GEN_2378; // @[Rob.scala 310:156 Rob.scala 310:156]
  wire [31:0] _GEN_2380 = 3'h4 == io_rob_init_info_bits_1_op1_rob ? rob_info_4_commit_data : _GEN_2379; // @[Rob.scala 310:156 Rob.scala 310:156]
  wire [31:0] _GEN_2381 = 3'h5 == io_rob_init_info_bits_1_op1_rob ? rob_info_5_commit_data : _GEN_2380; // @[Rob.scala 310:156 Rob.scala 310:156]
  wire [31:0] _GEN_2382 = 3'h6 == io_rob_init_info_bits_1_op1_rob ? rob_info_6_commit_data : _GEN_2381; // @[Rob.scala 310:156 Rob.scala 310:156]
  wire [31:0] _GEN_2383 = 3'h7 == io_rob_init_info_bits_1_op1_rob ? rob_info_7_commit_data : _GEN_2382; // @[Rob.scala 310:156 Rob.scala 310:156]
  wire  init_op1_hit_commit_1 = rob_commit_1_des_rob == io_rob_init_info_bits_1_op1_rob & rob_commit_valid_1 |
    rob_commit_0_des_rob == io_rob_init_info_bits_1_op1_rob & rob_commit_valid_0; // @[Rob.scala 359:92 Rob.scala 360:31]
  wire [31:0] _GEN_3481 = rob_commit_0_des_rob == io_rob_init_info_bits_1_op1_rob & rob_commit_valid_0 ?
    rob_commit_0_commit_data : 32'h0; // @[Rob.scala 359:92 Rob.scala 361:32]
  wire [31:0] init_op1_commit_data_1 = rob_commit_1_des_rob == io_rob_init_info_bits_1_op1_rob & rob_commit_valid_1 ?
    rob_commit_1_commit_data : _GEN_3481; // @[Rob.scala 359:92 Rob.scala 361:32]
  wire [31:0] _init_op1_data_T_4 = init_op1_hit_commit_1 ? init_op1_commit_data_1 : _GEN_2383; // @[Rob.scala 310:156]
  wire  init_op1_hit_wb_1 = io_wb_info_i_4_bits_rob_idx == io_rob_init_info_bits_1_op1_rob & io_wb_info_i_4_valid | (
    io_wb_info_i_3_bits_rob_idx == io_rob_init_info_bits_1_op1_rob & io_wb_info_i_3_valid | (io_wb_info_i_2_bits_rob_idx
     == io_rob_init_info_bits_1_op1_rob & io_wb_info_i_2_valid | (io_wb_info_i_1_bits_rob_idx ==
    io_rob_init_info_bits_1_op1_rob & io_wb_info_i_1_valid | io_wb_info_i_0_bits_rob_idx ==
    io_rob_init_info_bits_1_op1_rob & io_wb_info_i_0_valid))); // @[Rob.scala 371:101 Rob.scala 372:27]
  wire [31:0] _GEN_3509 = io_wb_info_i_0_bits_rob_idx == io_rob_init_info_bits_1_op1_rob & io_wb_info_i_0_valid ?
    io_wb_info_i_0_bits_data : 32'h0; // @[Rob.scala 371:101 Rob.scala 373:28]
  wire [31:0] _GEN_3513 = io_wb_info_i_1_bits_rob_idx == io_rob_init_info_bits_1_op1_rob & io_wb_info_i_1_valid ?
    io_wb_info_i_1_bits_data : _GEN_3509; // @[Rob.scala 371:101 Rob.scala 373:28]
  wire [31:0] _GEN_3517 = io_wb_info_i_2_bits_rob_idx == io_rob_init_info_bits_1_op1_rob & io_wb_info_i_2_valid ?
    io_wb_info_i_2_bits_data : _GEN_3513; // @[Rob.scala 371:101 Rob.scala 373:28]
  wire [31:0] _GEN_3521 = io_wb_info_i_3_bits_rob_idx == io_rob_init_info_bits_1_op1_rob & io_wb_info_i_3_valid ?
    io_wb_info_i_3_bits_data : _GEN_3517; // @[Rob.scala 371:101 Rob.scala 373:28]
  wire [31:0] init_op1_wb_data_1 = io_wb_info_i_4_bits_rob_idx == io_rob_init_info_bits_1_op1_rob & io_wb_info_i_4_valid
     ? io_wb_info_i_4_bits_data : _GEN_3521; // @[Rob.scala 371:101 Rob.scala 373:28]
  wire [31:0] _init_op1_data_T_5 = init_op1_hit_wb_1 ? init_op1_wb_data_1 : _init_op1_data_T_4; // @[Rob.scala 310:111]
  wire [31:0] init_op1_data_1 = ~io_rob_init_info_bits_1_op1_in_rob ? io_rob_init_info_bits_1_op1_regData :
    _init_op1_data_T_5; // @[Rob.scala 310:31]
  wire  _init_op2_data_T_3 = ~io_rob_init_info_bits_1_op2_in_rob; // @[Rob.scala 311:32]
  wire [31:0] _GEN_2385 = 3'h1 == io_rob_init_info_bits_1_op2_rob ? rob_info_1_commit_data : rob_info_0_commit_data; // @[Rob.scala 311:156 Rob.scala 311:156]
  wire [31:0] _GEN_2386 = 3'h2 == io_rob_init_info_bits_1_op2_rob ? rob_info_2_commit_data : _GEN_2385; // @[Rob.scala 311:156 Rob.scala 311:156]
  wire [31:0] _GEN_2387 = 3'h3 == io_rob_init_info_bits_1_op2_rob ? rob_info_3_commit_data : _GEN_2386; // @[Rob.scala 311:156 Rob.scala 311:156]
  wire [31:0] _GEN_2388 = 3'h4 == io_rob_init_info_bits_1_op2_rob ? rob_info_4_commit_data : _GEN_2387; // @[Rob.scala 311:156 Rob.scala 311:156]
  wire [31:0] _GEN_2389 = 3'h5 == io_rob_init_info_bits_1_op2_rob ? rob_info_5_commit_data : _GEN_2388; // @[Rob.scala 311:156 Rob.scala 311:156]
  wire [31:0] _GEN_2390 = 3'h6 == io_rob_init_info_bits_1_op2_rob ? rob_info_6_commit_data : _GEN_2389; // @[Rob.scala 311:156 Rob.scala 311:156]
  wire [31:0] _GEN_2391 = 3'h7 == io_rob_init_info_bits_1_op2_rob ? rob_info_7_commit_data : _GEN_2390; // @[Rob.scala 311:156 Rob.scala 311:156]
  wire  init_op2_hit_commit_1 = rob_commit_1_des_rob == io_rob_init_info_bits_1_op2_rob & rob_commit_valid_1 |
    rob_commit_0_des_rob == io_rob_init_info_bits_1_op2_rob & rob_commit_valid_0; // @[Rob.scala 363:92 Rob.scala 364:31]
  wire [31:0] _GEN_3483 = rob_commit_0_des_rob == io_rob_init_info_bits_1_op2_rob & rob_commit_valid_0 ?
    rob_commit_0_commit_data : 32'h0; // @[Rob.scala 363:92 Rob.scala 365:32]
  wire [31:0] init_op2_commit_data_1 = rob_commit_1_des_rob == io_rob_init_info_bits_1_op2_rob & rob_commit_valid_1 ?
    rob_commit_1_commit_data : _GEN_3483; // @[Rob.scala 363:92 Rob.scala 365:32]
  wire [31:0] _init_op2_data_T_4 = init_op2_hit_commit_1 ? init_op2_commit_data_1 : _GEN_2391; // @[Rob.scala 311:156]
  wire  init_op2_hit_wb_1 = io_wb_info_i_4_bits_rob_idx == io_rob_init_info_bits_1_op2_rob & io_wb_info_i_4_valid | (
    io_wb_info_i_3_bits_rob_idx == io_rob_init_info_bits_1_op2_rob & io_wb_info_i_3_valid | (io_wb_info_i_2_bits_rob_idx
     == io_rob_init_info_bits_1_op2_rob & io_wb_info_i_2_valid | (io_wb_info_i_1_bits_rob_idx ==
    io_rob_init_info_bits_1_op2_rob & io_wb_info_i_1_valid | io_wb_info_i_0_bits_rob_idx ==
    io_rob_init_info_bits_1_op2_rob & io_wb_info_i_0_valid))); // @[Rob.scala 375:101 Rob.scala 376:27]
  wire [31:0] _GEN_3511 = io_wb_info_i_0_bits_rob_idx == io_rob_init_info_bits_1_op2_rob & io_wb_info_i_0_valid ?
    io_wb_info_i_0_bits_data : 32'h0; // @[Rob.scala 375:101 Rob.scala 377:28]
  wire [31:0] _GEN_3515 = io_wb_info_i_1_bits_rob_idx == io_rob_init_info_bits_1_op2_rob & io_wb_info_i_1_valid ?
    io_wb_info_i_1_bits_data : _GEN_3511; // @[Rob.scala 375:101 Rob.scala 377:28]
  wire [31:0] _GEN_3519 = io_wb_info_i_2_bits_rob_idx == io_rob_init_info_bits_1_op2_rob & io_wb_info_i_2_valid ?
    io_wb_info_i_2_bits_data : _GEN_3515; // @[Rob.scala 375:101 Rob.scala 377:28]
  wire [31:0] _GEN_3523 = io_wb_info_i_3_bits_rob_idx == io_rob_init_info_bits_1_op2_rob & io_wb_info_i_3_valid ?
    io_wb_info_i_3_bits_data : _GEN_3519; // @[Rob.scala 375:101 Rob.scala 377:28]
  wire [31:0] init_op2_wb_data_1 = io_wb_info_i_4_bits_rob_idx == io_rob_init_info_bits_1_op2_rob & io_wb_info_i_4_valid
     ? io_wb_info_i_4_bits_data : _GEN_3523; // @[Rob.scala 375:101 Rob.scala 377:28]
  wire [31:0] _init_op2_data_T_5 = init_op2_hit_wb_1 ? init_op2_wb_data_1 : _init_op2_data_T_4; // @[Rob.scala 311:111]
  wire [31:0] init_op2_data_1 = ~io_rob_init_info_bits_1_op2_in_rob ? io_rob_init_info_bits_1_op2_regData :
    _init_op2_data_T_5; // @[Rob.scala 311:31]
  wire  _GEN_2393 = 3'h1 == io_rob_init_info_bits_1_op1_rob ? rob_info_1_commit_ready : rob_info_0_commit_ready; // @[Rob.scala 312:59 Rob.scala 312:59]
  wire  _GEN_2394 = 3'h2 == io_rob_init_info_bits_1_op1_rob ? rob_info_2_commit_ready : _GEN_2393; // @[Rob.scala 312:59 Rob.scala 312:59]
  wire  _GEN_2395 = 3'h3 == io_rob_init_info_bits_1_op1_rob ? rob_info_3_commit_ready : _GEN_2394; // @[Rob.scala 312:59 Rob.scala 312:59]
  wire  _GEN_2396 = 3'h4 == io_rob_init_info_bits_1_op1_rob ? rob_info_4_commit_ready : _GEN_2395; // @[Rob.scala 312:59 Rob.scala 312:59]
  wire  _GEN_2397 = 3'h5 == io_rob_init_info_bits_1_op1_rob ? rob_info_5_commit_ready : _GEN_2396; // @[Rob.scala 312:59 Rob.scala 312:59]
  wire  _GEN_2398 = 3'h6 == io_rob_init_info_bits_1_op1_rob ? rob_info_6_commit_ready : _GEN_2397; // @[Rob.scala 312:59 Rob.scala 312:59]
  wire  _GEN_2399 = 3'h7 == io_rob_init_info_bits_1_op1_rob ? rob_info_7_commit_ready : _GEN_2398; // @[Rob.scala 312:59 Rob.scala 312:59]
  wire  _GEN_2401 = 3'h1 == io_rob_init_info_bits_1_op1_rob ? rob_info_1_is_valid : rob_info_0_is_valid; // @[Rob.scala 312:59 Rob.scala 312:59]
  wire  _GEN_2402 = 3'h2 == io_rob_init_info_bits_1_op1_rob ? rob_info_2_is_valid : _GEN_2401; // @[Rob.scala 312:59 Rob.scala 312:59]
  wire  _GEN_2403 = 3'h3 == io_rob_init_info_bits_1_op1_rob ? rob_info_3_is_valid : _GEN_2402; // @[Rob.scala 312:59 Rob.scala 312:59]
  wire  _GEN_2404 = 3'h4 == io_rob_init_info_bits_1_op1_rob ? rob_info_4_is_valid : _GEN_2403; // @[Rob.scala 312:59 Rob.scala 312:59]
  wire  _GEN_2405 = 3'h5 == io_rob_init_info_bits_1_op1_rob ? rob_info_5_is_valid : _GEN_2404; // @[Rob.scala 312:59 Rob.scala 312:59]
  wire  _GEN_2406 = 3'h6 == io_rob_init_info_bits_1_op1_rob ? rob_info_6_is_valid : _GEN_2405; // @[Rob.scala 312:59 Rob.scala 312:59]
  wire  _GEN_2407 = 3'h7 == io_rob_init_info_bits_1_op1_rob ? rob_info_7_is_valid : _GEN_2406; // @[Rob.scala 312:59 Rob.scala 312:59]
  wire  init_op1_hit_rob_1 = _GEN_2399 & _GEN_2407 | init_op1_hit_wb_1 | init_op1_hit_commit_1; // @[Rob.scala 312:111]
  wire  _GEN_2409 = 3'h1 == io_rob_init_info_bits_1_op2_rob ? rob_info_1_commit_ready : rob_info_0_commit_ready; // @[Rob.scala 313:59 Rob.scala 313:59]
  wire  _GEN_2410 = 3'h2 == io_rob_init_info_bits_1_op2_rob ? rob_info_2_commit_ready : _GEN_2409; // @[Rob.scala 313:59 Rob.scala 313:59]
  wire  _GEN_2411 = 3'h3 == io_rob_init_info_bits_1_op2_rob ? rob_info_3_commit_ready : _GEN_2410; // @[Rob.scala 313:59 Rob.scala 313:59]
  wire  _GEN_2412 = 3'h4 == io_rob_init_info_bits_1_op2_rob ? rob_info_4_commit_ready : _GEN_2411; // @[Rob.scala 313:59 Rob.scala 313:59]
  wire  _GEN_2413 = 3'h5 == io_rob_init_info_bits_1_op2_rob ? rob_info_5_commit_ready : _GEN_2412; // @[Rob.scala 313:59 Rob.scala 313:59]
  wire  _GEN_2414 = 3'h6 == io_rob_init_info_bits_1_op2_rob ? rob_info_6_commit_ready : _GEN_2413; // @[Rob.scala 313:59 Rob.scala 313:59]
  wire  _GEN_2415 = 3'h7 == io_rob_init_info_bits_1_op2_rob ? rob_info_7_commit_ready : _GEN_2414; // @[Rob.scala 313:59 Rob.scala 313:59]
  wire  _GEN_2417 = 3'h1 == io_rob_init_info_bits_1_op2_rob ? rob_info_1_is_valid : rob_info_0_is_valid; // @[Rob.scala 313:59 Rob.scala 313:59]
  wire  _GEN_2418 = 3'h2 == io_rob_init_info_bits_1_op2_rob ? rob_info_2_is_valid : _GEN_2417; // @[Rob.scala 313:59 Rob.scala 313:59]
  wire  _GEN_2419 = 3'h3 == io_rob_init_info_bits_1_op2_rob ? rob_info_3_is_valid : _GEN_2418; // @[Rob.scala 313:59 Rob.scala 313:59]
  wire  _GEN_2420 = 3'h4 == io_rob_init_info_bits_1_op2_rob ? rob_info_4_is_valid : _GEN_2419; // @[Rob.scala 313:59 Rob.scala 313:59]
  wire  _GEN_2421 = 3'h5 == io_rob_init_info_bits_1_op2_rob ? rob_info_5_is_valid : _GEN_2420; // @[Rob.scala 313:59 Rob.scala 313:59]
  wire  _GEN_2422 = 3'h6 == io_rob_init_info_bits_1_op2_rob ? rob_info_6_is_valid : _GEN_2421; // @[Rob.scala 313:59 Rob.scala 313:59]
  wire  _GEN_2423 = 3'h7 == io_rob_init_info_bits_1_op2_rob ? rob_info_7_is_valid : _GEN_2422; // @[Rob.scala 313:59 Rob.scala 313:59]
  wire  init_op2_hit_rob_1 = _GEN_2415 & _GEN_2423 | init_op2_hit_wb_1 | init_op2_hit_commit_1; // @[Rob.scala 313:111]
  wire [31:0] _GEN_2424 = 3'h0 == io_rob_init_info_bits_1_des_rob ? init_op1_data_1 : _GEN_2320; // @[Rob.scala 316:34 Rob.scala 316:34]
  wire [31:0] _GEN_2425 = 3'h1 == io_rob_init_info_bits_1_des_rob ? init_op1_data_1 : _GEN_2321; // @[Rob.scala 316:34 Rob.scala 316:34]
  wire [31:0] _GEN_2426 = 3'h2 == io_rob_init_info_bits_1_des_rob ? init_op1_data_1 : _GEN_2322; // @[Rob.scala 316:34 Rob.scala 316:34]
  wire [31:0] _GEN_2427 = 3'h3 == io_rob_init_info_bits_1_des_rob ? init_op1_data_1 : _GEN_2323; // @[Rob.scala 316:34 Rob.scala 316:34]
  wire [31:0] _GEN_2428 = 3'h4 == io_rob_init_info_bits_1_des_rob ? init_op1_data_1 : _GEN_2324; // @[Rob.scala 316:34 Rob.scala 316:34]
  wire [31:0] _GEN_2429 = 3'h5 == io_rob_init_info_bits_1_des_rob ? init_op1_data_1 : _GEN_2325; // @[Rob.scala 316:34 Rob.scala 316:34]
  wire [31:0] _GEN_2430 = 3'h6 == io_rob_init_info_bits_1_des_rob ? init_op1_data_1 : _GEN_2326; // @[Rob.scala 316:34 Rob.scala 316:34]
  wire [31:0] _GEN_2431 = 3'h7 == io_rob_init_info_bits_1_des_rob ? init_op1_data_1 : _GEN_2327; // @[Rob.scala 316:34 Rob.scala 316:34]
  wire [31:0] _GEN_2432 = 3'h0 == io_rob_init_info_bits_1_des_rob ? init_op2_data_1 : _GEN_2328; // @[Rob.scala 317:34 Rob.scala 317:34]
  wire [31:0] _GEN_2433 = 3'h1 == io_rob_init_info_bits_1_des_rob ? init_op2_data_1 : _GEN_2329; // @[Rob.scala 317:34 Rob.scala 317:34]
  wire [31:0] _GEN_2434 = 3'h2 == io_rob_init_info_bits_1_des_rob ? init_op2_data_1 : _GEN_2330; // @[Rob.scala 317:34 Rob.scala 317:34]
  wire [31:0] _GEN_2435 = 3'h3 == io_rob_init_info_bits_1_des_rob ? init_op2_data_1 : _GEN_2331; // @[Rob.scala 317:34 Rob.scala 317:34]
  wire [31:0] _GEN_2436 = 3'h4 == io_rob_init_info_bits_1_des_rob ? init_op2_data_1 : _GEN_2332; // @[Rob.scala 317:34 Rob.scala 317:34]
  wire [31:0] _GEN_2437 = 3'h5 == io_rob_init_info_bits_1_des_rob ? init_op2_data_1 : _GEN_2333; // @[Rob.scala 317:34 Rob.scala 317:34]
  wire [31:0] _GEN_2438 = 3'h6 == io_rob_init_info_bits_1_des_rob ? init_op2_data_1 : _GEN_2334; // @[Rob.scala 317:34 Rob.scala 317:34]
  wire [31:0] _GEN_2439 = 3'h7 == io_rob_init_info_bits_1_des_rob ? init_op2_data_1 : _GEN_2335; // @[Rob.scala 317:34 Rob.scala 317:34]
  wire [2:0] _GEN_2440 = 3'h0 == io_rob_init_info_bits_1_des_rob ? io_rob_init_info_bits_1_op1_rob : _GEN_2336; // @[Rob.scala 318:33 Rob.scala 318:33]
  wire [2:0] _GEN_2441 = 3'h1 == io_rob_init_info_bits_1_des_rob ? io_rob_init_info_bits_1_op1_rob : _GEN_2337; // @[Rob.scala 318:33 Rob.scala 318:33]
  wire [2:0] _GEN_2442 = 3'h2 == io_rob_init_info_bits_1_des_rob ? io_rob_init_info_bits_1_op1_rob : _GEN_2338; // @[Rob.scala 318:33 Rob.scala 318:33]
  wire [2:0] _GEN_2443 = 3'h3 == io_rob_init_info_bits_1_des_rob ? io_rob_init_info_bits_1_op1_rob : _GEN_2339; // @[Rob.scala 318:33 Rob.scala 318:33]
  wire [2:0] _GEN_2444 = 3'h4 == io_rob_init_info_bits_1_des_rob ? io_rob_init_info_bits_1_op1_rob : _GEN_2340; // @[Rob.scala 318:33 Rob.scala 318:33]
  wire [2:0] _GEN_2445 = 3'h5 == io_rob_init_info_bits_1_des_rob ? io_rob_init_info_bits_1_op1_rob : _GEN_2341; // @[Rob.scala 318:33 Rob.scala 318:33]
  wire [2:0] _GEN_2446 = 3'h6 == io_rob_init_info_bits_1_des_rob ? io_rob_init_info_bits_1_op1_rob : _GEN_2342; // @[Rob.scala 318:33 Rob.scala 318:33]
  wire [2:0] _GEN_2447 = 3'h7 == io_rob_init_info_bits_1_des_rob ? io_rob_init_info_bits_1_op1_rob : _GEN_2343; // @[Rob.scala 318:33 Rob.scala 318:33]
  wire [2:0] _GEN_2448 = 3'h0 == io_rob_init_info_bits_1_des_rob ? io_rob_init_info_bits_1_op2_rob : _GEN_2344; // @[Rob.scala 319:33 Rob.scala 319:33]
  wire [2:0] _GEN_2449 = 3'h1 == io_rob_init_info_bits_1_des_rob ? io_rob_init_info_bits_1_op2_rob : _GEN_2345; // @[Rob.scala 319:33 Rob.scala 319:33]
  wire [2:0] _GEN_2450 = 3'h2 == io_rob_init_info_bits_1_des_rob ? io_rob_init_info_bits_1_op2_rob : _GEN_2346; // @[Rob.scala 319:33 Rob.scala 319:33]
  wire [2:0] _GEN_2451 = 3'h3 == io_rob_init_info_bits_1_des_rob ? io_rob_init_info_bits_1_op2_rob : _GEN_2347; // @[Rob.scala 319:33 Rob.scala 319:33]
  wire [2:0] _GEN_2452 = 3'h4 == io_rob_init_info_bits_1_des_rob ? io_rob_init_info_bits_1_op2_rob : _GEN_2348; // @[Rob.scala 319:33 Rob.scala 319:33]
  wire [2:0] _GEN_2453 = 3'h5 == io_rob_init_info_bits_1_des_rob ? io_rob_init_info_bits_1_op2_rob : _GEN_2349; // @[Rob.scala 319:33 Rob.scala 319:33]
  wire [2:0] _GEN_2454 = 3'h6 == io_rob_init_info_bits_1_des_rob ? io_rob_init_info_bits_1_op2_rob : _GEN_2350; // @[Rob.scala 319:33 Rob.scala 319:33]
  wire [2:0] _GEN_2455 = 3'h7 == io_rob_init_info_bits_1_des_rob ? io_rob_init_info_bits_1_op2_rob : _GEN_2351; // @[Rob.scala 319:33 Rob.scala 319:33]
  wire  _GEN_2456 = 3'h0 == io_rob_init_info_bits_1_des_rob ? _init_op1_data_T_3 | init_op1_hit_rob_1 : _GEN_2352; // @[Rob.scala 320:35 Rob.scala 320:35]
  wire  _GEN_2457 = 3'h1 == io_rob_init_info_bits_1_des_rob ? _init_op1_data_T_3 | init_op1_hit_rob_1 : _GEN_2353; // @[Rob.scala 320:35 Rob.scala 320:35]
  wire  _GEN_2458 = 3'h2 == io_rob_init_info_bits_1_des_rob ? _init_op1_data_T_3 | init_op1_hit_rob_1 : _GEN_2354; // @[Rob.scala 320:35 Rob.scala 320:35]
  wire  _GEN_2459 = 3'h3 == io_rob_init_info_bits_1_des_rob ? _init_op1_data_T_3 | init_op1_hit_rob_1 : _GEN_2355; // @[Rob.scala 320:35 Rob.scala 320:35]
  wire  _GEN_2460 = 3'h4 == io_rob_init_info_bits_1_des_rob ? _init_op1_data_T_3 | init_op1_hit_rob_1 : _GEN_2356; // @[Rob.scala 320:35 Rob.scala 320:35]
  wire  _GEN_2461 = 3'h5 == io_rob_init_info_bits_1_des_rob ? _init_op1_data_T_3 | init_op1_hit_rob_1 : _GEN_2357; // @[Rob.scala 320:35 Rob.scala 320:35]
  wire  _GEN_2462 = 3'h6 == io_rob_init_info_bits_1_des_rob ? _init_op1_data_T_3 | init_op1_hit_rob_1 : _GEN_2358; // @[Rob.scala 320:35 Rob.scala 320:35]
  wire  _GEN_2463 = 3'h7 == io_rob_init_info_bits_1_des_rob ? _init_op1_data_T_3 | init_op1_hit_rob_1 : _GEN_2359; // @[Rob.scala 320:35 Rob.scala 320:35]
  wire  _GEN_2464 = 3'h0 == io_rob_init_info_bits_1_des_rob ? _init_op2_data_T_3 | init_op2_hit_rob_1 : _GEN_2360; // @[Rob.scala 321:35 Rob.scala 321:35]
  wire  _GEN_2465 = 3'h1 == io_rob_init_info_bits_1_des_rob ? _init_op2_data_T_3 | init_op2_hit_rob_1 : _GEN_2361; // @[Rob.scala 321:35 Rob.scala 321:35]
  wire  _GEN_2466 = 3'h2 == io_rob_init_info_bits_1_des_rob ? _init_op2_data_T_3 | init_op2_hit_rob_1 : _GEN_2362; // @[Rob.scala 321:35 Rob.scala 321:35]
  wire  _GEN_2467 = 3'h3 == io_rob_init_info_bits_1_des_rob ? _init_op2_data_T_3 | init_op2_hit_rob_1 : _GEN_2363; // @[Rob.scala 321:35 Rob.scala 321:35]
  wire  _GEN_2468 = 3'h4 == io_rob_init_info_bits_1_des_rob ? _init_op2_data_T_3 | init_op2_hit_rob_1 : _GEN_2364; // @[Rob.scala 321:35 Rob.scala 321:35]
  wire  _GEN_2469 = 3'h5 == io_rob_init_info_bits_1_des_rob ? _init_op2_data_T_3 | init_op2_hit_rob_1 : _GEN_2365; // @[Rob.scala 321:35 Rob.scala 321:35]
  wire  _GEN_2470 = 3'h6 == io_rob_init_info_bits_1_des_rob ? _init_op2_data_T_3 | init_op2_hit_rob_1 : _GEN_2366; // @[Rob.scala 321:35 Rob.scala 321:35]
  wire  _GEN_2471 = 3'h7 == io_rob_init_info_bits_1_des_rob ? _init_op2_data_T_3 | init_op2_hit_rob_1 : _GEN_2367; // @[Rob.scala 321:35 Rob.scala 321:35]
  wire  _GEN_2472 = 3'h0 == io_rob_init_info_bits_1_des_rob | _GEN_2368; // @[Rob.scala 322:33 Rob.scala 322:33]
  wire  _GEN_2473 = 3'h1 == io_rob_init_info_bits_1_des_rob | _GEN_2369; // @[Rob.scala 322:33 Rob.scala 322:33]
  wire  _GEN_2474 = 3'h2 == io_rob_init_info_bits_1_des_rob | _GEN_2370; // @[Rob.scala 322:33 Rob.scala 322:33]
  wire  _GEN_2475 = 3'h3 == io_rob_init_info_bits_1_des_rob | _GEN_2371; // @[Rob.scala 322:33 Rob.scala 322:33]
  wire  _GEN_2476 = 3'h4 == io_rob_init_info_bits_1_des_rob | _GEN_2372; // @[Rob.scala 322:33 Rob.scala 322:33]
  wire  _GEN_2477 = 3'h5 == io_rob_init_info_bits_1_des_rob | _GEN_2373; // @[Rob.scala 322:33 Rob.scala 322:33]
  wire  _GEN_2478 = 3'h6 == io_rob_init_info_bits_1_des_rob | _GEN_2374; // @[Rob.scala 322:33 Rob.scala 322:33]
  wire  _GEN_2479 = 3'h7 == io_rob_init_info_bits_1_des_rob | _GEN_2375; // @[Rob.scala 322:33 Rob.scala 322:33]
  wire [31:0] _GEN_2480 = io_rob_init_info_valid & io_rob_init_info_bits_1_is_valid & _T_21 ? _GEN_2424 : _GEN_2320; // @[Rob.scala 315:86]
  wire [31:0] _GEN_2481 = io_rob_init_info_valid & io_rob_init_info_bits_1_is_valid & _T_21 ? _GEN_2425 : _GEN_2321; // @[Rob.scala 315:86]
  wire [31:0] _GEN_2482 = io_rob_init_info_valid & io_rob_init_info_bits_1_is_valid & _T_21 ? _GEN_2426 : _GEN_2322; // @[Rob.scala 315:86]
  wire [31:0] _GEN_2483 = io_rob_init_info_valid & io_rob_init_info_bits_1_is_valid & _T_21 ? _GEN_2427 : _GEN_2323; // @[Rob.scala 315:86]
  wire [31:0] _GEN_2484 = io_rob_init_info_valid & io_rob_init_info_bits_1_is_valid & _T_21 ? _GEN_2428 : _GEN_2324; // @[Rob.scala 315:86]
  wire [31:0] _GEN_2485 = io_rob_init_info_valid & io_rob_init_info_bits_1_is_valid & _T_21 ? _GEN_2429 : _GEN_2325; // @[Rob.scala 315:86]
  wire [31:0] _GEN_2486 = io_rob_init_info_valid & io_rob_init_info_bits_1_is_valid & _T_21 ? _GEN_2430 : _GEN_2326; // @[Rob.scala 315:86]
  wire [31:0] _GEN_2487 = io_rob_init_info_valid & io_rob_init_info_bits_1_is_valid & _T_21 ? _GEN_2431 : _GEN_2327; // @[Rob.scala 315:86]
  wire [31:0] _GEN_2488 = io_rob_init_info_valid & io_rob_init_info_bits_1_is_valid & _T_21 ? _GEN_2432 : _GEN_2328; // @[Rob.scala 315:86]
  wire [31:0] _GEN_2489 = io_rob_init_info_valid & io_rob_init_info_bits_1_is_valid & _T_21 ? _GEN_2433 : _GEN_2329; // @[Rob.scala 315:86]
  wire [31:0] _GEN_2490 = io_rob_init_info_valid & io_rob_init_info_bits_1_is_valid & _T_21 ? _GEN_2434 : _GEN_2330; // @[Rob.scala 315:86]
  wire [31:0] _GEN_2491 = io_rob_init_info_valid & io_rob_init_info_bits_1_is_valid & _T_21 ? _GEN_2435 : _GEN_2331; // @[Rob.scala 315:86]
  wire [31:0] _GEN_2492 = io_rob_init_info_valid & io_rob_init_info_bits_1_is_valid & _T_21 ? _GEN_2436 : _GEN_2332; // @[Rob.scala 315:86]
  wire [31:0] _GEN_2493 = io_rob_init_info_valid & io_rob_init_info_bits_1_is_valid & _T_21 ? _GEN_2437 : _GEN_2333; // @[Rob.scala 315:86]
  wire [31:0] _GEN_2494 = io_rob_init_info_valid & io_rob_init_info_bits_1_is_valid & _T_21 ? _GEN_2438 : _GEN_2334; // @[Rob.scala 315:86]
  wire [31:0] _GEN_2495 = io_rob_init_info_valid & io_rob_init_info_bits_1_is_valid & _T_21 ? _GEN_2439 : _GEN_2335; // @[Rob.scala 315:86]
  wire [2:0] _GEN_2496 = io_rob_init_info_valid & io_rob_init_info_bits_1_is_valid & _T_21 ? _GEN_2440 : _GEN_2336; // @[Rob.scala 315:86]
  wire [2:0] _GEN_2497 = io_rob_init_info_valid & io_rob_init_info_bits_1_is_valid & _T_21 ? _GEN_2441 : _GEN_2337; // @[Rob.scala 315:86]
  wire [2:0] _GEN_2498 = io_rob_init_info_valid & io_rob_init_info_bits_1_is_valid & _T_21 ? _GEN_2442 : _GEN_2338; // @[Rob.scala 315:86]
  wire [2:0] _GEN_2499 = io_rob_init_info_valid & io_rob_init_info_bits_1_is_valid & _T_21 ? _GEN_2443 : _GEN_2339; // @[Rob.scala 315:86]
  wire [2:0] _GEN_2500 = io_rob_init_info_valid & io_rob_init_info_bits_1_is_valid & _T_21 ? _GEN_2444 : _GEN_2340; // @[Rob.scala 315:86]
  wire [2:0] _GEN_2501 = io_rob_init_info_valid & io_rob_init_info_bits_1_is_valid & _T_21 ? _GEN_2445 : _GEN_2341; // @[Rob.scala 315:86]
  wire [2:0] _GEN_2502 = io_rob_init_info_valid & io_rob_init_info_bits_1_is_valid & _T_21 ? _GEN_2446 : _GEN_2342; // @[Rob.scala 315:86]
  wire [2:0] _GEN_2503 = io_rob_init_info_valid & io_rob_init_info_bits_1_is_valid & _T_21 ? _GEN_2447 : _GEN_2343; // @[Rob.scala 315:86]
  wire [2:0] _GEN_2504 = io_rob_init_info_valid & io_rob_init_info_bits_1_is_valid & _T_21 ? _GEN_2448 : _GEN_2344; // @[Rob.scala 315:86]
  wire [2:0] _GEN_2505 = io_rob_init_info_valid & io_rob_init_info_bits_1_is_valid & _T_21 ? _GEN_2449 : _GEN_2345; // @[Rob.scala 315:86]
  wire [2:0] _GEN_2506 = io_rob_init_info_valid & io_rob_init_info_bits_1_is_valid & _T_21 ? _GEN_2450 : _GEN_2346; // @[Rob.scala 315:86]
  wire [2:0] _GEN_2507 = io_rob_init_info_valid & io_rob_init_info_bits_1_is_valid & _T_21 ? _GEN_2451 : _GEN_2347; // @[Rob.scala 315:86]
  wire [2:0] _GEN_2508 = io_rob_init_info_valid & io_rob_init_info_bits_1_is_valid & _T_21 ? _GEN_2452 : _GEN_2348; // @[Rob.scala 315:86]
  wire [2:0] _GEN_2509 = io_rob_init_info_valid & io_rob_init_info_bits_1_is_valid & _T_21 ? _GEN_2453 : _GEN_2349; // @[Rob.scala 315:86]
  wire [2:0] _GEN_2510 = io_rob_init_info_valid & io_rob_init_info_bits_1_is_valid & _T_21 ? _GEN_2454 : _GEN_2350; // @[Rob.scala 315:86]
  wire [2:0] _GEN_2511 = io_rob_init_info_valid & io_rob_init_info_bits_1_is_valid & _T_21 ? _GEN_2455 : _GEN_2351; // @[Rob.scala 315:86]
  wire  _GEN_2512 = io_rob_init_info_valid & io_rob_init_info_bits_1_is_valid & _T_21 ? _GEN_2456 : _GEN_2352; // @[Rob.scala 315:86]
  wire  _GEN_2513 = io_rob_init_info_valid & io_rob_init_info_bits_1_is_valid & _T_21 ? _GEN_2457 : _GEN_2353; // @[Rob.scala 315:86]
  wire  _GEN_2514 = io_rob_init_info_valid & io_rob_init_info_bits_1_is_valid & _T_21 ? _GEN_2458 : _GEN_2354; // @[Rob.scala 315:86]
  wire  _GEN_2515 = io_rob_init_info_valid & io_rob_init_info_bits_1_is_valid & _T_21 ? _GEN_2459 : _GEN_2355; // @[Rob.scala 315:86]
  wire  _GEN_2516 = io_rob_init_info_valid & io_rob_init_info_bits_1_is_valid & _T_21 ? _GEN_2460 : _GEN_2356; // @[Rob.scala 315:86]
  wire  _GEN_2517 = io_rob_init_info_valid & io_rob_init_info_bits_1_is_valid & _T_21 ? _GEN_2461 : _GEN_2357; // @[Rob.scala 315:86]
  wire  _GEN_2518 = io_rob_init_info_valid & io_rob_init_info_bits_1_is_valid & _T_21 ? _GEN_2462 : _GEN_2358; // @[Rob.scala 315:86]
  wire  _GEN_2519 = io_rob_init_info_valid & io_rob_init_info_bits_1_is_valid & _T_21 ? _GEN_2463 : _GEN_2359; // @[Rob.scala 315:86]
  wire  _GEN_2520 = io_rob_init_info_valid & io_rob_init_info_bits_1_is_valid & _T_21 ? _GEN_2464 : _GEN_2360; // @[Rob.scala 315:86]
  wire  _GEN_2521 = io_rob_init_info_valid & io_rob_init_info_bits_1_is_valid & _T_21 ? _GEN_2465 : _GEN_2361; // @[Rob.scala 315:86]
  wire  _GEN_2522 = io_rob_init_info_valid & io_rob_init_info_bits_1_is_valid & _T_21 ? _GEN_2466 : _GEN_2362; // @[Rob.scala 315:86]
  wire  _GEN_2523 = io_rob_init_info_valid & io_rob_init_info_bits_1_is_valid & _T_21 ? _GEN_2467 : _GEN_2363; // @[Rob.scala 315:86]
  wire  _GEN_2524 = io_rob_init_info_valid & io_rob_init_info_bits_1_is_valid & _T_21 ? _GEN_2468 : _GEN_2364; // @[Rob.scala 315:86]
  wire  _GEN_2525 = io_rob_init_info_valid & io_rob_init_info_bits_1_is_valid & _T_21 ? _GEN_2469 : _GEN_2365; // @[Rob.scala 315:86]
  wire  _GEN_2526 = io_rob_init_info_valid & io_rob_init_info_bits_1_is_valid & _T_21 ? _GEN_2470 : _GEN_2366; // @[Rob.scala 315:86]
  wire  _GEN_2527 = io_rob_init_info_valid & io_rob_init_info_bits_1_is_valid & _T_21 ? _GEN_2471 : _GEN_2367; // @[Rob.scala 315:86]
  wire  _GEN_2528 = io_rob_init_info_valid & io_rob_init_info_bits_1_is_valid & _T_21 ? _GEN_2472 : _GEN_2368; // @[Rob.scala 315:86]
  wire  _GEN_2529 = io_rob_init_info_valid & io_rob_init_info_bits_1_is_valid & _T_21 ? _GEN_2473 : _GEN_2369; // @[Rob.scala 315:86]
  wire  _GEN_2530 = io_rob_init_info_valid & io_rob_init_info_bits_1_is_valid & _T_21 ? _GEN_2474 : _GEN_2370; // @[Rob.scala 315:86]
  wire  _GEN_2531 = io_rob_init_info_valid & io_rob_init_info_bits_1_is_valid & _T_21 ? _GEN_2475 : _GEN_2371; // @[Rob.scala 315:86]
  wire  _GEN_2532 = io_rob_init_info_valid & io_rob_init_info_bits_1_is_valid & _T_21 ? _GEN_2476 : _GEN_2372; // @[Rob.scala 315:86]
  wire  _GEN_2533 = io_rob_init_info_valid & io_rob_init_info_bits_1_is_valid & _T_21 ? _GEN_2477 : _GEN_2373; // @[Rob.scala 315:86]
  wire  _GEN_2534 = io_rob_init_info_valid & io_rob_init_info_bits_1_is_valid & _T_21 ? _GEN_2478 : _GEN_2374; // @[Rob.scala 315:86]
  wire  _GEN_2535 = io_rob_init_info_valid & io_rob_init_info_bits_1_is_valid & _T_21 ? _GEN_2479 : _GEN_2375; // @[Rob.scala 315:86]
  wire  commit_ready_mask_0 = _GEN_7 & _GEN_23; // @[Rob.scala 329:67]
  wire  commit_ready_mask_1 = _GEN_47 & _GEN_63; // @[Rob.scala 329:67]
  wire  commit_wait_mask_0 = ~commit_ready_mask_0; // @[Rob.scala 330:48]
  wire  commit_wait_mask_1 = ~commit_ready_mask_1; // @[Rob.scala 330:48]
  wire  _GEN_2569 = 3'h1 == dispatch_idxs_0 ? rob_info_1_predict_miss : rob_info_0_predict_miss; // @[Rob.scala 331:73 Rob.scala 331:73]
  wire  _GEN_2570 = 3'h2 == dispatch_idxs_0 ? rob_info_2_predict_miss : _GEN_2569; // @[Rob.scala 331:73 Rob.scala 331:73]
  wire  _GEN_2571 = 3'h3 == dispatch_idxs_0 ? rob_info_3_predict_miss : _GEN_2570; // @[Rob.scala 331:73 Rob.scala 331:73]
  wire  _GEN_2572 = 3'h4 == dispatch_idxs_0 ? rob_info_4_predict_miss : _GEN_2571; // @[Rob.scala 331:73 Rob.scala 331:73]
  wire  _GEN_2573 = 3'h5 == dispatch_idxs_0 ? rob_info_5_predict_miss : _GEN_2572; // @[Rob.scala 331:73 Rob.scala 331:73]
  wire  _GEN_2574 = 3'h6 == dispatch_idxs_0 ? rob_info_6_predict_miss : _GEN_2573; // @[Rob.scala 331:73 Rob.scala 331:73]
  wire  _GEN_2575 = 3'h7 == dispatch_idxs_0 ? rob_info_7_predict_miss : _GEN_2574; // @[Rob.scala 331:73 Rob.scala 331:73]
  wire  _GEN_2577 = 3'h1 == dispatch_idxs_0 ? rob_info_1_flush_on_commit : rob_info_0_flush_on_commit; // @[Rob.scala 331:73 Rob.scala 331:73]
  wire  _GEN_2578 = 3'h2 == dispatch_idxs_0 ? rob_info_2_flush_on_commit : _GEN_2577; // @[Rob.scala 331:73 Rob.scala 331:73]
  wire  _GEN_2579 = 3'h3 == dispatch_idxs_0 ? rob_info_3_flush_on_commit : _GEN_2578; // @[Rob.scala 331:73 Rob.scala 331:73]
  wire  _GEN_2580 = 3'h4 == dispatch_idxs_0 ? rob_info_4_flush_on_commit : _GEN_2579; // @[Rob.scala 331:73 Rob.scala 331:73]
  wire  _GEN_2581 = 3'h5 == dispatch_idxs_0 ? rob_info_5_flush_on_commit : _GEN_2580; // @[Rob.scala 331:73 Rob.scala 331:73]
  wire  _GEN_2582 = 3'h6 == dispatch_idxs_0 ? rob_info_6_flush_on_commit : _GEN_2581; // @[Rob.scala 331:73 Rob.scala 331:73]
  wire  _GEN_2583 = 3'h7 == dispatch_idxs_0 ? rob_info_7_flush_on_commit : _GEN_2582; // @[Rob.scala 331:73 Rob.scala 331:73]
  wire  need_flush_mask_0 = _GEN_2575 | _GEN_2583; // @[Rob.scala 331:73]
  wire  _GEN_2585 = 3'h1 == dispatch_idxs_1 ? rob_info_1_predict_miss : rob_info_0_predict_miss; // @[Rob.scala 331:73 Rob.scala 331:73]
  wire  _GEN_2586 = 3'h2 == dispatch_idxs_1 ? rob_info_2_predict_miss : _GEN_2585; // @[Rob.scala 331:73 Rob.scala 331:73]
  wire  _GEN_2587 = 3'h3 == dispatch_idxs_1 ? rob_info_3_predict_miss : _GEN_2586; // @[Rob.scala 331:73 Rob.scala 331:73]
  wire  _GEN_2588 = 3'h4 == dispatch_idxs_1 ? rob_info_4_predict_miss : _GEN_2587; // @[Rob.scala 331:73 Rob.scala 331:73]
  wire  _GEN_2589 = 3'h5 == dispatch_idxs_1 ? rob_info_5_predict_miss : _GEN_2588; // @[Rob.scala 331:73 Rob.scala 331:73]
  wire  _GEN_2590 = 3'h6 == dispatch_idxs_1 ? rob_info_6_predict_miss : _GEN_2589; // @[Rob.scala 331:73 Rob.scala 331:73]
  wire  _GEN_2591 = 3'h7 == dispatch_idxs_1 ? rob_info_7_predict_miss : _GEN_2590; // @[Rob.scala 331:73 Rob.scala 331:73]
  wire  _GEN_2593 = 3'h1 == dispatch_idxs_1 ? rob_info_1_flush_on_commit : rob_info_0_flush_on_commit; // @[Rob.scala 331:73 Rob.scala 331:73]
  wire  _GEN_2594 = 3'h2 == dispatch_idxs_1 ? rob_info_2_flush_on_commit : _GEN_2593; // @[Rob.scala 331:73 Rob.scala 331:73]
  wire  _GEN_2595 = 3'h3 == dispatch_idxs_1 ? rob_info_3_flush_on_commit : _GEN_2594; // @[Rob.scala 331:73 Rob.scala 331:73]
  wire  _GEN_2596 = 3'h4 == dispatch_idxs_1 ? rob_info_4_flush_on_commit : _GEN_2595; // @[Rob.scala 331:73 Rob.scala 331:73]
  wire  _GEN_2597 = 3'h5 == dispatch_idxs_1 ? rob_info_5_flush_on_commit : _GEN_2596; // @[Rob.scala 331:73 Rob.scala 331:73]
  wire  _GEN_2598 = 3'h6 == dispatch_idxs_1 ? rob_info_6_flush_on_commit : _GEN_2597; // @[Rob.scala 331:73 Rob.scala 331:73]
  wire  _GEN_2599 = 3'h7 == dispatch_idxs_1 ? rob_info_7_flush_on_commit : _GEN_2598; // @[Rob.scala 331:73 Rob.scala 331:73]
  wire  need_flush_mask_1 = _GEN_2591 | _GEN_2599; // @[Rob.scala 331:73]
  wire  deq_wait_mask_1 = commit_wait_mask_0 | need_flush_mask_0 | commit_wait_mask_1; // @[Rob.scala 332:133]
  wire [1:0] _head_next_T = deq_wait_mask_1 ? 2'h1 : 2'h2; // @[Mux.scala 47:69]
  wire [1:0] _head_next_T_1 = commit_wait_mask_0 ? 2'h0 : _head_next_T; // @[Mux.scala 47:69]
  wire  deq_ready_mask_0 = ~commit_wait_mask_0; // @[Rob.scala 334:50]
  wire  deq_ready_mask_1 = ~deq_wait_mask_1; // @[Rob.scala 334:50]
  wire  flush_idx = need_flush_mask_0 ? 1'h0 : 1'h1; // @[Mux.scala 47:69]
  wire  _GEN_2604 = flush_idx ? need_flush_mask_1 : need_flush_mask_0; // @[Rob.scala 337:52 Rob.scala 337:52]
  wire  _GEN_2606 = flush_idx ? deq_ready_mask_1 : deq_ready_mask_0; // @[Rob.scala 337:52 Rob.scala 337:52]
  wire [1:0] _GEN_4151 = {{1'd0}, flush_idx}; // @[Rob.scala 337:52 Rob.scala 337:52]
  wire  flush = _GEN_2604 & (2'h2 == _GEN_4151 | _GEN_2606); // @[Rob.scala 337:52]
  reg [4:0] rob_commit_0_commit_addr; // @[Rob.scala 341:23]
  reg [4:0] rob_commit_1_commit_addr; // @[Rob.scala 341:23]
  wire [31:0] _GEN_2609 = 3'h1 == dispatch_idxs_0 ? rob_info_1_commit_data : rob_info_0_commit_data; // @[Rob.scala 346:31 Rob.scala 346:31]
  wire [31:0] _GEN_2610 = 3'h2 == dispatch_idxs_0 ? rob_info_2_commit_data : _GEN_2609; // @[Rob.scala 346:31 Rob.scala 346:31]
  wire [31:0] _GEN_2611 = 3'h3 == dispatch_idxs_0 ? rob_info_3_commit_data : _GEN_2610; // @[Rob.scala 346:31 Rob.scala 346:31]
  wire [31:0] _GEN_2612 = 3'h4 == dispatch_idxs_0 ? rob_info_4_commit_data : _GEN_2611; // @[Rob.scala 346:31 Rob.scala 346:31]
  wire [31:0] _GEN_2613 = 3'h5 == dispatch_idxs_0 ? rob_info_5_commit_data : _GEN_2612; // @[Rob.scala 346:31 Rob.scala 346:31]
  wire [4:0] _GEN_2617 = 3'h1 == dispatch_idxs_0 ? rob_info_1_commit_addr : rob_info_0_commit_addr; // @[Rob.scala 348:31 Rob.scala 348:31]
  wire [4:0] _GEN_2618 = 3'h2 == dispatch_idxs_0 ? rob_info_2_commit_addr : _GEN_2617; // @[Rob.scala 348:31 Rob.scala 348:31]
  wire [4:0] _GEN_2619 = 3'h3 == dispatch_idxs_0 ? rob_info_3_commit_addr : _GEN_2618; // @[Rob.scala 348:31 Rob.scala 348:31]
  wire [4:0] _GEN_2620 = 3'h4 == dispatch_idxs_0 ? rob_info_4_commit_addr : _GEN_2619; // @[Rob.scala 348:31 Rob.scala 348:31]
  wire [4:0] _GEN_2621 = 3'h5 == dispatch_idxs_0 ? rob_info_5_commit_addr : _GEN_2620; // @[Rob.scala 348:31 Rob.scala 348:31]
  wire  _GEN_2624 = 3'h0 == dispatch_idxs_0 ? 1'h0 : _GEN_1384; // @[Rob.scala 42:13 Rob.scala 42:13]
  wire  _GEN_2625 = 3'h1 == dispatch_idxs_0 ? 1'h0 : _GEN_1385; // @[Rob.scala 42:13 Rob.scala 42:13]
  wire  _GEN_2626 = 3'h2 == dispatch_idxs_0 ? 1'h0 : _GEN_1386; // @[Rob.scala 42:13 Rob.scala 42:13]
  wire  _GEN_2627 = 3'h3 == dispatch_idxs_0 ? 1'h0 : _GEN_1387; // @[Rob.scala 42:13 Rob.scala 42:13]
  wire  _GEN_2628 = 3'h4 == dispatch_idxs_0 ? 1'h0 : _GEN_1388; // @[Rob.scala 42:13 Rob.scala 42:13]
  wire  _GEN_2629 = 3'h5 == dispatch_idxs_0 ? 1'h0 : _GEN_1389; // @[Rob.scala 42:13 Rob.scala 42:13]
  wire  _GEN_2630 = 3'h6 == dispatch_idxs_0 ? 1'h0 : _GEN_1390; // @[Rob.scala 42:13 Rob.scala 42:13]
  wire  _GEN_2631 = 3'h7 == dispatch_idxs_0 ? 1'h0 : _GEN_1391; // @[Rob.scala 42:13 Rob.scala 42:13]
  wire  _GEN_2632 = 3'h0 == dispatch_idxs_0 ? 1'h0 : _GEN_2184; // @[Rob.scala 43:9 Rob.scala 43:9]
  wire  _GEN_2633 = 3'h1 == dispatch_idxs_0 ? 1'h0 : _GEN_2185; // @[Rob.scala 43:9 Rob.scala 43:9]
  wire  _GEN_2634 = 3'h2 == dispatch_idxs_0 ? 1'h0 : _GEN_2186; // @[Rob.scala 43:9 Rob.scala 43:9]
  wire  _GEN_2635 = 3'h3 == dispatch_idxs_0 ? 1'h0 : _GEN_2187; // @[Rob.scala 43:9 Rob.scala 43:9]
  wire  _GEN_2636 = 3'h4 == dispatch_idxs_0 ? 1'h0 : _GEN_2188; // @[Rob.scala 43:9 Rob.scala 43:9]
  wire  _GEN_2637 = 3'h5 == dispatch_idxs_0 ? 1'h0 : _GEN_2189; // @[Rob.scala 43:9 Rob.scala 43:9]
  wire  _GEN_2638 = 3'h6 == dispatch_idxs_0 ? 1'h0 : _GEN_2190; // @[Rob.scala 43:9 Rob.scala 43:9]
  wire  _GEN_2639 = 3'h7 == dispatch_idxs_0 ? 1'h0 : _GEN_2191; // @[Rob.scala 43:9 Rob.scala 43:9]
  wire [5:0] _GEN_2640 = 3'h0 == dispatch_idxs_0 ? 6'h0 : _GEN_1488; // @[Rob.scala 44:8 Rob.scala 44:8]
  wire [5:0] _GEN_2641 = 3'h1 == dispatch_idxs_0 ? 6'h0 : _GEN_1489; // @[Rob.scala 44:8 Rob.scala 44:8]
  wire [5:0] _GEN_2642 = 3'h2 == dispatch_idxs_0 ? 6'h0 : _GEN_1490; // @[Rob.scala 44:8 Rob.scala 44:8]
  wire [5:0] _GEN_2643 = 3'h3 == dispatch_idxs_0 ? 6'h0 : _GEN_1491; // @[Rob.scala 44:8 Rob.scala 44:8]
  wire [5:0] _GEN_2644 = 3'h4 == dispatch_idxs_0 ? 6'h0 : _GEN_1492; // @[Rob.scala 44:8 Rob.scala 44:8]
  wire [5:0] _GEN_2645 = 3'h5 == dispatch_idxs_0 ? 6'h0 : _GEN_1493; // @[Rob.scala 44:8 Rob.scala 44:8]
  wire [5:0] _GEN_2646 = 3'h6 == dispatch_idxs_0 ? 6'h0 : _GEN_1494; // @[Rob.scala 44:8 Rob.scala 44:8]
  wire [5:0] _GEN_2647 = 3'h7 == dispatch_idxs_0 ? 6'h0 : _GEN_1495; // @[Rob.scala 44:8 Rob.scala 44:8]
  wire [2:0] _GEN_2648 = 3'h0 == dispatch_idxs_0 ? 3'h0 : _GEN_1496; // @[Rob.scala 45:13 Rob.scala 45:13]
  wire [2:0] _GEN_2649 = 3'h1 == dispatch_idxs_0 ? 3'h0 : _GEN_1497; // @[Rob.scala 45:13 Rob.scala 45:13]
  wire [2:0] _GEN_2650 = 3'h2 == dispatch_idxs_0 ? 3'h0 : _GEN_1498; // @[Rob.scala 45:13 Rob.scala 45:13]
  wire [2:0] _GEN_2651 = 3'h3 == dispatch_idxs_0 ? 3'h0 : _GEN_1499; // @[Rob.scala 45:13 Rob.scala 45:13]
  wire [2:0] _GEN_2652 = 3'h4 == dispatch_idxs_0 ? 3'h0 : _GEN_1500; // @[Rob.scala 45:13 Rob.scala 45:13]
  wire [2:0] _GEN_2653 = 3'h5 == dispatch_idxs_0 ? 3'h0 : _GEN_1501; // @[Rob.scala 45:13 Rob.scala 45:13]
  wire [2:0] _GEN_2654 = 3'h6 == dispatch_idxs_0 ? 3'h0 : _GEN_1502; // @[Rob.scala 45:13 Rob.scala 45:13]
  wire [2:0] _GEN_2655 = 3'h7 == dispatch_idxs_0 ? 3'h0 : _GEN_1503; // @[Rob.scala 45:13 Rob.scala 45:13]
  wire  _GEN_2656 = 3'h0 == dispatch_idxs_0 ? 1'h0 : _GEN_1504; // @[Rob.scala 46:13 Rob.scala 46:13]
  wire  _GEN_2657 = 3'h1 == dispatch_idxs_0 ? 1'h0 : _GEN_1505; // @[Rob.scala 46:13 Rob.scala 46:13]
  wire  _GEN_2658 = 3'h2 == dispatch_idxs_0 ? 1'h0 : _GEN_1506; // @[Rob.scala 46:13 Rob.scala 46:13]
  wire  _GEN_2659 = 3'h3 == dispatch_idxs_0 ? 1'h0 : _GEN_1507; // @[Rob.scala 46:13 Rob.scala 46:13]
  wire  _GEN_2660 = 3'h4 == dispatch_idxs_0 ? 1'h0 : _GEN_1508; // @[Rob.scala 46:13 Rob.scala 46:13]
  wire  _GEN_2661 = 3'h5 == dispatch_idxs_0 ? 1'h0 : _GEN_1509; // @[Rob.scala 46:13 Rob.scala 46:13]
  wire  _GEN_2662 = 3'h6 == dispatch_idxs_0 ? 1'h0 : _GEN_1510; // @[Rob.scala 46:13 Rob.scala 46:13]
  wire  _GEN_2663 = 3'h7 == dispatch_idxs_0 ? 1'h0 : _GEN_1511; // @[Rob.scala 46:13 Rob.scala 46:13]
  wire [31:0] _GEN_2664 = 3'h0 == dispatch_idxs_0 ? 32'h0 : _GEN_1432; // @[Rob.scala 47:14 Rob.scala 47:14]
  wire [31:0] _GEN_2665 = 3'h1 == dispatch_idxs_0 ? 32'h0 : _GEN_1433; // @[Rob.scala 47:14 Rob.scala 47:14]
  wire [31:0] _GEN_2666 = 3'h2 == dispatch_idxs_0 ? 32'h0 : _GEN_1434; // @[Rob.scala 47:14 Rob.scala 47:14]
  wire [31:0] _GEN_2667 = 3'h3 == dispatch_idxs_0 ? 32'h0 : _GEN_1435; // @[Rob.scala 47:14 Rob.scala 47:14]
  wire [31:0] _GEN_2668 = 3'h4 == dispatch_idxs_0 ? 32'h0 : _GEN_1436; // @[Rob.scala 47:14 Rob.scala 47:14]
  wire [31:0] _GEN_2669 = 3'h5 == dispatch_idxs_0 ? 32'h0 : _GEN_1437; // @[Rob.scala 47:14 Rob.scala 47:14]
  wire [31:0] _GEN_2670 = 3'h6 == dispatch_idxs_0 ? 32'h0 : _GEN_1438; // @[Rob.scala 47:14 Rob.scala 47:14]
  wire [31:0] _GEN_2671 = 3'h7 == dispatch_idxs_0 ? 32'h0 : _GEN_1439; // @[Rob.scala 47:14 Rob.scala 47:14]
  wire [4:0] _GEN_2672 = 3'h0 == dispatch_idxs_0 ? 5'h0 : _GEN_1440; // @[Rob.scala 48:16 Rob.scala 48:16]
  wire [4:0] _GEN_2673 = 3'h1 == dispatch_idxs_0 ? 5'h0 : _GEN_1441; // @[Rob.scala 48:16 Rob.scala 48:16]
  wire [4:0] _GEN_2674 = 3'h2 == dispatch_idxs_0 ? 5'h0 : _GEN_1442; // @[Rob.scala 48:16 Rob.scala 48:16]
  wire [4:0] _GEN_2675 = 3'h3 == dispatch_idxs_0 ? 5'h0 : _GEN_1443; // @[Rob.scala 48:16 Rob.scala 48:16]
  wire [4:0] _GEN_2676 = 3'h4 == dispatch_idxs_0 ? 5'h0 : _GEN_1444; // @[Rob.scala 48:16 Rob.scala 48:16]
  wire [4:0] _GEN_2677 = 3'h5 == dispatch_idxs_0 ? 5'h0 : _GEN_1445; // @[Rob.scala 48:16 Rob.scala 48:16]
  wire [4:0] _GEN_2678 = 3'h6 == dispatch_idxs_0 ? 5'h0 : _GEN_1446; // @[Rob.scala 48:16 Rob.scala 48:16]
  wire [4:0] _GEN_2679 = 3'h7 == dispatch_idxs_0 ? 5'h0 : _GEN_1447; // @[Rob.scala 48:16 Rob.scala 48:16]
  wire [31:0] _GEN_2680 = 3'h0 == dispatch_idxs_0 ? 32'h0 : _GEN_2168; // @[Rob.scala 49:16 Rob.scala 49:16]
  wire [31:0] _GEN_2681 = 3'h1 == dispatch_idxs_0 ? 32'h0 : _GEN_2169; // @[Rob.scala 49:16 Rob.scala 49:16]
  wire [31:0] _GEN_2682 = 3'h2 == dispatch_idxs_0 ? 32'h0 : _GEN_2170; // @[Rob.scala 49:16 Rob.scala 49:16]
  wire [31:0] _GEN_2683 = 3'h3 == dispatch_idxs_0 ? 32'h0 : _GEN_2171; // @[Rob.scala 49:16 Rob.scala 49:16]
  wire [31:0] _GEN_2684 = 3'h4 == dispatch_idxs_0 ? 32'h0 : _GEN_2172; // @[Rob.scala 49:16 Rob.scala 49:16]
  wire [31:0] _GEN_2685 = 3'h5 == dispatch_idxs_0 ? 32'h0 : _GEN_2173; // @[Rob.scala 49:16 Rob.scala 49:16]
  wire [31:0] _GEN_2686 = 3'h6 == dispatch_idxs_0 ? 32'h0 : _GEN_2174; // @[Rob.scala 49:16 Rob.scala 49:16]
  wire [31:0] _GEN_2687 = 3'h7 == dispatch_idxs_0 ? 32'h0 : _GEN_2175; // @[Rob.scala 49:16 Rob.scala 49:16]
  wire  _GEN_2696 = 3'h0 == dispatch_idxs_0 ? 1'h0 : _GEN_2176; // @[Rob.scala 51:17 Rob.scala 51:17]
  wire  _GEN_2697 = 3'h1 == dispatch_idxs_0 ? 1'h0 : _GEN_2177; // @[Rob.scala 51:17 Rob.scala 51:17]
  wire  _GEN_2698 = 3'h2 == dispatch_idxs_0 ? 1'h0 : _GEN_2178; // @[Rob.scala 51:17 Rob.scala 51:17]
  wire  _GEN_2699 = 3'h3 == dispatch_idxs_0 ? 1'h0 : _GEN_2179; // @[Rob.scala 51:17 Rob.scala 51:17]
  wire  _GEN_2700 = 3'h4 == dispatch_idxs_0 ? 1'h0 : _GEN_2180; // @[Rob.scala 51:17 Rob.scala 51:17]
  wire  _GEN_2701 = 3'h5 == dispatch_idxs_0 ? 1'h0 : _GEN_2181; // @[Rob.scala 51:17 Rob.scala 51:17]
  wire  _GEN_2702 = 3'h6 == dispatch_idxs_0 ? 1'h0 : _GEN_2182; // @[Rob.scala 51:17 Rob.scala 51:17]
  wire  _GEN_2703 = 3'h7 == dispatch_idxs_0 ? 1'h0 : _GEN_2183; // @[Rob.scala 51:17 Rob.scala 51:17]
  wire  _GEN_2712 = 3'h0 == dispatch_idxs_0 ? 1'h0 : _GEN_1464; // @[Rob.scala 53:14 Rob.scala 53:14]
  wire  _GEN_2713 = 3'h1 == dispatch_idxs_0 ? 1'h0 : _GEN_1465; // @[Rob.scala 53:14 Rob.scala 53:14]
  wire  _GEN_2714 = 3'h2 == dispatch_idxs_0 ? 1'h0 : _GEN_1466; // @[Rob.scala 53:14 Rob.scala 53:14]
  wire  _GEN_2715 = 3'h3 == dispatch_idxs_0 ? 1'h0 : _GEN_1467; // @[Rob.scala 53:14 Rob.scala 53:14]
  wire  _GEN_2716 = 3'h4 == dispatch_idxs_0 ? 1'h0 : _GEN_1468; // @[Rob.scala 53:14 Rob.scala 53:14]
  wire  _GEN_2717 = 3'h5 == dispatch_idxs_0 ? 1'h0 : _GEN_1469; // @[Rob.scala 53:14 Rob.scala 53:14]
  wire  _GEN_2718 = 3'h6 == dispatch_idxs_0 ? 1'h0 : _GEN_1470; // @[Rob.scala 53:14 Rob.scala 53:14]
  wire  _GEN_2719 = 3'h7 == dispatch_idxs_0 ? 1'h0 : _GEN_1471; // @[Rob.scala 53:14 Rob.scala 53:14]
  wire  _GEN_2728 = 3'h0 == dispatch_idxs_0 ? 1'h0 : _GEN_1528; // @[Rob.scala 55:18 Rob.scala 55:18]
  wire  _GEN_2729 = 3'h1 == dispatch_idxs_0 ? 1'h0 : _GEN_1529; // @[Rob.scala 55:18 Rob.scala 55:18]
  wire  _GEN_2730 = 3'h2 == dispatch_idxs_0 ? 1'h0 : _GEN_1530; // @[Rob.scala 55:18 Rob.scala 55:18]
  wire  _GEN_2731 = 3'h3 == dispatch_idxs_0 ? 1'h0 : _GEN_1531; // @[Rob.scala 55:18 Rob.scala 55:18]
  wire  _GEN_2732 = 3'h4 == dispatch_idxs_0 ? 1'h0 : _GEN_1532; // @[Rob.scala 55:18 Rob.scala 55:18]
  wire  _GEN_2733 = 3'h5 == dispatch_idxs_0 ? 1'h0 : _GEN_1533; // @[Rob.scala 55:18 Rob.scala 55:18]
  wire  _GEN_2734 = 3'h6 == dispatch_idxs_0 ? 1'h0 : _GEN_1534; // @[Rob.scala 55:18 Rob.scala 55:18]
  wire  _GEN_2735 = 3'h7 == dispatch_idxs_0 ? 1'h0 : _GEN_1535; // @[Rob.scala 55:18 Rob.scala 55:18]
  wire  _GEN_2736 = 3'h0 == dispatch_idxs_0 ? 1'h0 : _GEN_2192; // @[Rob.scala 56:13 Rob.scala 56:13]
  wire  _GEN_2737 = 3'h1 == dispatch_idxs_0 ? 1'h0 : _GEN_2193; // @[Rob.scala 56:13 Rob.scala 56:13]
  wire  _GEN_2738 = 3'h2 == dispatch_idxs_0 ? 1'h0 : _GEN_2194; // @[Rob.scala 56:13 Rob.scala 56:13]
  wire  _GEN_2739 = 3'h3 == dispatch_idxs_0 ? 1'h0 : _GEN_2195; // @[Rob.scala 56:13 Rob.scala 56:13]
  wire  _GEN_2740 = 3'h4 == dispatch_idxs_0 ? 1'h0 : _GEN_2196; // @[Rob.scala 56:13 Rob.scala 56:13]
  wire  _GEN_2741 = 3'h5 == dispatch_idxs_0 ? 1'h0 : _GEN_2197; // @[Rob.scala 56:13 Rob.scala 56:13]
  wire  _GEN_2742 = 3'h6 == dispatch_idxs_0 ? 1'h0 : _GEN_2198; // @[Rob.scala 56:13 Rob.scala 56:13]
  wire  _GEN_2743 = 3'h7 == dispatch_idxs_0 ? 1'h0 : _GEN_2199; // @[Rob.scala 56:13 Rob.scala 56:13]
  wire  _GEN_2744 = 3'h0 == dispatch_idxs_0 ? 1'h0 : _GEN_2200; // @[Rob.scala 57:17 Rob.scala 57:17]
  wire  _GEN_2745 = 3'h1 == dispatch_idxs_0 ? 1'h0 : _GEN_2201; // @[Rob.scala 57:17 Rob.scala 57:17]
  wire  _GEN_2746 = 3'h2 == dispatch_idxs_0 ? 1'h0 : _GEN_2202; // @[Rob.scala 57:17 Rob.scala 57:17]
  wire  _GEN_2747 = 3'h3 == dispatch_idxs_0 ? 1'h0 : _GEN_2203; // @[Rob.scala 57:17 Rob.scala 57:17]
  wire  _GEN_2748 = 3'h4 == dispatch_idxs_0 ? 1'h0 : _GEN_2204; // @[Rob.scala 57:17 Rob.scala 57:17]
  wire  _GEN_2749 = 3'h5 == dispatch_idxs_0 ? 1'h0 : _GEN_2205; // @[Rob.scala 57:17 Rob.scala 57:17]
  wire  _GEN_2750 = 3'h6 == dispatch_idxs_0 ? 1'h0 : _GEN_2206; // @[Rob.scala 57:17 Rob.scala 57:17]
  wire  _GEN_2751 = 3'h7 == dispatch_idxs_0 ? 1'h0 : _GEN_2207; // @[Rob.scala 57:17 Rob.scala 57:17]
  wire [3:0] _GEN_2752 = 3'h0 == dispatch_idxs_0 ? 4'h0 : _GEN_1480; // @[Rob.scala 58:12 Rob.scala 58:12]
  wire [3:0] _GEN_2753 = 3'h1 == dispatch_idxs_0 ? 4'h0 : _GEN_1481; // @[Rob.scala 58:12 Rob.scala 58:12]
  wire [3:0] _GEN_2754 = 3'h2 == dispatch_idxs_0 ? 4'h0 : _GEN_1482; // @[Rob.scala 58:12 Rob.scala 58:12]
  wire [3:0] _GEN_2755 = 3'h3 == dispatch_idxs_0 ? 4'h0 : _GEN_1483; // @[Rob.scala 58:12 Rob.scala 58:12]
  wire [3:0] _GEN_2756 = 3'h4 == dispatch_idxs_0 ? 4'h0 : _GEN_1484; // @[Rob.scala 58:12 Rob.scala 58:12]
  wire [3:0] _GEN_2757 = 3'h5 == dispatch_idxs_0 ? 4'h0 : _GEN_1485; // @[Rob.scala 58:12 Rob.scala 58:12]
  wire [3:0] _GEN_2758 = 3'h6 == dispatch_idxs_0 ? 4'h0 : _GEN_1486; // @[Rob.scala 58:12 Rob.scala 58:12]
  wire [3:0] _GEN_2759 = 3'h7 == dispatch_idxs_0 ? 4'h0 : _GEN_1487; // @[Rob.scala 58:12 Rob.scala 58:12]
  wire  _GEN_2760 = 3'h0 == dispatch_idxs_0 ? 1'h0 : _GEN_2512; // @[Rob.scala 59:14 Rob.scala 59:14]
  wire  _GEN_2761 = 3'h1 == dispatch_idxs_0 ? 1'h0 : _GEN_2513; // @[Rob.scala 59:14 Rob.scala 59:14]
  wire  _GEN_2762 = 3'h2 == dispatch_idxs_0 ? 1'h0 : _GEN_2514; // @[Rob.scala 59:14 Rob.scala 59:14]
  wire  _GEN_2763 = 3'h3 == dispatch_idxs_0 ? 1'h0 : _GEN_2515; // @[Rob.scala 59:14 Rob.scala 59:14]
  wire  _GEN_2764 = 3'h4 == dispatch_idxs_0 ? 1'h0 : _GEN_2516; // @[Rob.scala 59:14 Rob.scala 59:14]
  wire  _GEN_2765 = 3'h5 == dispatch_idxs_0 ? 1'h0 : _GEN_2517; // @[Rob.scala 59:14 Rob.scala 59:14]
  wire  _GEN_2766 = 3'h6 == dispatch_idxs_0 ? 1'h0 : _GEN_2518; // @[Rob.scala 59:14 Rob.scala 59:14]
  wire  _GEN_2767 = 3'h7 == dispatch_idxs_0 ? 1'h0 : _GEN_2519; // @[Rob.scala 59:14 Rob.scala 59:14]
  wire [2:0] _GEN_2768 = 3'h0 == dispatch_idxs_0 ? 3'h0 : _GEN_2496; // @[Rob.scala 60:12 Rob.scala 60:12]
  wire [2:0] _GEN_2769 = 3'h1 == dispatch_idxs_0 ? 3'h0 : _GEN_2497; // @[Rob.scala 60:12 Rob.scala 60:12]
  wire [2:0] _GEN_2770 = 3'h2 == dispatch_idxs_0 ? 3'h0 : _GEN_2498; // @[Rob.scala 60:12 Rob.scala 60:12]
  wire [2:0] _GEN_2771 = 3'h3 == dispatch_idxs_0 ? 3'h0 : _GEN_2499; // @[Rob.scala 60:12 Rob.scala 60:12]
  wire [2:0] _GEN_2772 = 3'h4 == dispatch_idxs_0 ? 3'h0 : _GEN_2500; // @[Rob.scala 60:12 Rob.scala 60:12]
  wire [2:0] _GEN_2773 = 3'h5 == dispatch_idxs_0 ? 3'h0 : _GEN_2501; // @[Rob.scala 60:12 Rob.scala 60:12]
  wire [2:0] _GEN_2774 = 3'h6 == dispatch_idxs_0 ? 3'h0 : _GEN_2502; // @[Rob.scala 60:12 Rob.scala 60:12]
  wire [2:0] _GEN_2775 = 3'h7 == dispatch_idxs_0 ? 3'h0 : _GEN_2503; // @[Rob.scala 60:12 Rob.scala 60:12]
  wire [31:0] _GEN_2776 = 3'h0 == dispatch_idxs_0 ? 32'h0 : _GEN_2480; // @[Rob.scala 61:13 Rob.scala 61:13]
  wire [31:0] _GEN_2777 = 3'h1 == dispatch_idxs_0 ? 32'h0 : _GEN_2481; // @[Rob.scala 61:13 Rob.scala 61:13]
  wire [31:0] _GEN_2778 = 3'h2 == dispatch_idxs_0 ? 32'h0 : _GEN_2482; // @[Rob.scala 61:13 Rob.scala 61:13]
  wire [31:0] _GEN_2779 = 3'h3 == dispatch_idxs_0 ? 32'h0 : _GEN_2483; // @[Rob.scala 61:13 Rob.scala 61:13]
  wire [31:0] _GEN_2780 = 3'h4 == dispatch_idxs_0 ? 32'h0 : _GEN_2484; // @[Rob.scala 61:13 Rob.scala 61:13]
  wire [31:0] _GEN_2781 = 3'h5 == dispatch_idxs_0 ? 32'h0 : _GEN_2485; // @[Rob.scala 61:13 Rob.scala 61:13]
  wire [31:0] _GEN_2782 = 3'h6 == dispatch_idxs_0 ? 32'h0 : _GEN_2486; // @[Rob.scala 61:13 Rob.scala 61:13]
  wire [31:0] _GEN_2783 = 3'h7 == dispatch_idxs_0 ? 32'h0 : _GEN_2487; // @[Rob.scala 61:13 Rob.scala 61:13]
  wire  _GEN_2784 = 3'h0 == dispatch_idxs_0 ? 1'h0 : _GEN_2520; // @[Rob.scala 62:14 Rob.scala 62:14]
  wire  _GEN_2785 = 3'h1 == dispatch_idxs_0 ? 1'h0 : _GEN_2521; // @[Rob.scala 62:14 Rob.scala 62:14]
  wire  _GEN_2786 = 3'h2 == dispatch_idxs_0 ? 1'h0 : _GEN_2522; // @[Rob.scala 62:14 Rob.scala 62:14]
  wire  _GEN_2787 = 3'h3 == dispatch_idxs_0 ? 1'h0 : _GEN_2523; // @[Rob.scala 62:14 Rob.scala 62:14]
  wire  _GEN_2788 = 3'h4 == dispatch_idxs_0 ? 1'h0 : _GEN_2524; // @[Rob.scala 62:14 Rob.scala 62:14]
  wire  _GEN_2789 = 3'h5 == dispatch_idxs_0 ? 1'h0 : _GEN_2525; // @[Rob.scala 62:14 Rob.scala 62:14]
  wire  _GEN_2790 = 3'h6 == dispatch_idxs_0 ? 1'h0 : _GEN_2526; // @[Rob.scala 62:14 Rob.scala 62:14]
  wire  _GEN_2791 = 3'h7 == dispatch_idxs_0 ? 1'h0 : _GEN_2527; // @[Rob.scala 62:14 Rob.scala 62:14]
  wire [2:0] _GEN_2792 = 3'h0 == dispatch_idxs_0 ? 3'h0 : _GEN_2504; // @[Rob.scala 63:12 Rob.scala 63:12]
  wire [2:0] _GEN_2793 = 3'h1 == dispatch_idxs_0 ? 3'h0 : _GEN_2505; // @[Rob.scala 63:12 Rob.scala 63:12]
  wire [2:0] _GEN_2794 = 3'h2 == dispatch_idxs_0 ? 3'h0 : _GEN_2506; // @[Rob.scala 63:12 Rob.scala 63:12]
  wire [2:0] _GEN_2795 = 3'h3 == dispatch_idxs_0 ? 3'h0 : _GEN_2507; // @[Rob.scala 63:12 Rob.scala 63:12]
  wire [2:0] _GEN_2796 = 3'h4 == dispatch_idxs_0 ? 3'h0 : _GEN_2508; // @[Rob.scala 63:12 Rob.scala 63:12]
  wire [2:0] _GEN_2797 = 3'h5 == dispatch_idxs_0 ? 3'h0 : _GEN_2509; // @[Rob.scala 63:12 Rob.scala 63:12]
  wire [2:0] _GEN_2798 = 3'h6 == dispatch_idxs_0 ? 3'h0 : _GEN_2510; // @[Rob.scala 63:12 Rob.scala 63:12]
  wire [2:0] _GEN_2799 = 3'h7 == dispatch_idxs_0 ? 3'h0 : _GEN_2511; // @[Rob.scala 63:12 Rob.scala 63:12]
  wire [31:0] _GEN_2800 = 3'h0 == dispatch_idxs_0 ? 32'h0 : _GEN_2488; // @[Rob.scala 64:13 Rob.scala 64:13]
  wire [31:0] _GEN_2801 = 3'h1 == dispatch_idxs_0 ? 32'h0 : _GEN_2489; // @[Rob.scala 64:13 Rob.scala 64:13]
  wire [31:0] _GEN_2802 = 3'h2 == dispatch_idxs_0 ? 32'h0 : _GEN_2490; // @[Rob.scala 64:13 Rob.scala 64:13]
  wire [31:0] _GEN_2803 = 3'h3 == dispatch_idxs_0 ? 32'h0 : _GEN_2491; // @[Rob.scala 64:13 Rob.scala 64:13]
  wire [31:0] _GEN_2804 = 3'h4 == dispatch_idxs_0 ? 32'h0 : _GEN_2492; // @[Rob.scala 64:13 Rob.scala 64:13]
  wire [31:0] _GEN_2805 = 3'h5 == dispatch_idxs_0 ? 32'h0 : _GEN_2493; // @[Rob.scala 64:13 Rob.scala 64:13]
  wire [31:0] _GEN_2806 = 3'h6 == dispatch_idxs_0 ? 32'h0 : _GEN_2494; // @[Rob.scala 64:13 Rob.scala 64:13]
  wire [31:0] _GEN_2807 = 3'h7 == dispatch_idxs_0 ? 32'h0 : _GEN_2495; // @[Rob.scala 64:13 Rob.scala 64:13]
  wire [31:0] _GEN_2808 = 3'h0 == dispatch_idxs_0 ? 32'h0 : _GEN_2208; // @[Rob.scala 65:13 Rob.scala 65:13]
  wire [31:0] _GEN_2809 = 3'h1 == dispatch_idxs_0 ? 32'h0 : _GEN_2209; // @[Rob.scala 65:13 Rob.scala 65:13]
  wire [31:0] _GEN_2810 = 3'h2 == dispatch_idxs_0 ? 32'h0 : _GEN_2210; // @[Rob.scala 65:13 Rob.scala 65:13]
  wire [31:0] _GEN_2811 = 3'h3 == dispatch_idxs_0 ? 32'h0 : _GEN_2211; // @[Rob.scala 65:13 Rob.scala 65:13]
  wire [31:0] _GEN_2812 = 3'h4 == dispatch_idxs_0 ? 32'h0 : _GEN_2212; // @[Rob.scala 65:13 Rob.scala 65:13]
  wire [31:0] _GEN_2813 = 3'h5 == dispatch_idxs_0 ? 32'h0 : _GEN_2213; // @[Rob.scala 65:13 Rob.scala 65:13]
  wire [31:0] _GEN_2814 = 3'h6 == dispatch_idxs_0 ? 32'h0 : _GEN_2214; // @[Rob.scala 65:13 Rob.scala 65:13]
  wire [31:0] _GEN_2815 = 3'h7 == dispatch_idxs_0 ? 32'h0 : _GEN_2215; // @[Rob.scala 65:13 Rob.scala 65:13]
  wire  _GEN_2816 = 3'h0 == dispatch_idxs_0 ? 1'h0 : _GEN_2528; // @[Rob.scala 66:13 Rob.scala 66:13]
  wire  _GEN_2817 = 3'h1 == dispatch_idxs_0 ? 1'h0 : _GEN_2529; // @[Rob.scala 66:13 Rob.scala 66:13]
  wire  _GEN_2818 = 3'h2 == dispatch_idxs_0 ? 1'h0 : _GEN_2530; // @[Rob.scala 66:13 Rob.scala 66:13]
  wire  _GEN_2819 = 3'h3 == dispatch_idxs_0 ? 1'h0 : _GEN_2531; // @[Rob.scala 66:13 Rob.scala 66:13]
  wire  _GEN_2820 = 3'h4 == dispatch_idxs_0 ? 1'h0 : _GEN_2532; // @[Rob.scala 66:13 Rob.scala 66:13]
  wire  _GEN_2821 = 3'h5 == dispatch_idxs_0 ? 1'h0 : _GEN_2533; // @[Rob.scala 66:13 Rob.scala 66:13]
  wire  _GEN_2822 = 3'h6 == dispatch_idxs_0 ? 1'h0 : _GEN_2534; // @[Rob.scala 66:13 Rob.scala 66:13]
  wire  _GEN_2823 = 3'h7 == dispatch_idxs_0 ? 1'h0 : _GEN_2535; // @[Rob.scala 66:13 Rob.scala 66:13]
  wire  _GEN_2824 = 3'h0 == dispatch_idxs_0 ? 1'h0 : _GEN_1520; // @[Rob.scala 67:20 Rob.scala 67:20]
  wire  _GEN_2825 = 3'h1 == dispatch_idxs_0 ? 1'h0 : _GEN_1521; // @[Rob.scala 67:20 Rob.scala 67:20]
  wire  _GEN_2826 = 3'h2 == dispatch_idxs_0 ? 1'h0 : _GEN_1522; // @[Rob.scala 67:20 Rob.scala 67:20]
  wire  _GEN_2827 = 3'h3 == dispatch_idxs_0 ? 1'h0 : _GEN_1523; // @[Rob.scala 67:20 Rob.scala 67:20]
  wire  _GEN_2828 = 3'h4 == dispatch_idxs_0 ? 1'h0 : _GEN_1524; // @[Rob.scala 67:20 Rob.scala 67:20]
  wire  _GEN_2829 = 3'h5 == dispatch_idxs_0 ? 1'h0 : _GEN_1525; // @[Rob.scala 67:20 Rob.scala 67:20]
  wire  _GEN_2830 = 3'h6 == dispatch_idxs_0 ? 1'h0 : _GEN_1526; // @[Rob.scala 67:20 Rob.scala 67:20]
  wire  _GEN_2831 = 3'h7 == dispatch_idxs_0 ? 1'h0 : _GEN_1527; // @[Rob.scala 67:20 Rob.scala 67:20]
  wire  _GEN_2832 = deq_ready_mask_0 ? _GEN_2624 : _GEN_1384; // @[Rob.scala 349:28]
  wire  _GEN_2833 = deq_ready_mask_0 ? _GEN_2625 : _GEN_1385; // @[Rob.scala 349:28]
  wire  _GEN_2834 = deq_ready_mask_0 ? _GEN_2626 : _GEN_1386; // @[Rob.scala 349:28]
  wire  _GEN_2835 = deq_ready_mask_0 ? _GEN_2627 : _GEN_1387; // @[Rob.scala 349:28]
  wire  _GEN_2836 = deq_ready_mask_0 ? _GEN_2628 : _GEN_1388; // @[Rob.scala 349:28]
  wire  _GEN_2837 = deq_ready_mask_0 ? _GEN_2629 : _GEN_1389; // @[Rob.scala 349:28]
  wire  _GEN_2838 = deq_ready_mask_0 ? _GEN_2630 : _GEN_1390; // @[Rob.scala 349:28]
  wire  _GEN_2839 = deq_ready_mask_0 ? _GEN_2631 : _GEN_1391; // @[Rob.scala 349:28]
  wire  _GEN_2840 = deq_ready_mask_0 ? _GEN_2632 : _GEN_2184; // @[Rob.scala 349:28]
  wire  _GEN_2841 = deq_ready_mask_0 ? _GEN_2633 : _GEN_2185; // @[Rob.scala 349:28]
  wire  _GEN_2842 = deq_ready_mask_0 ? _GEN_2634 : _GEN_2186; // @[Rob.scala 349:28]
  wire  _GEN_2843 = deq_ready_mask_0 ? _GEN_2635 : _GEN_2187; // @[Rob.scala 349:28]
  wire  _GEN_2844 = deq_ready_mask_0 ? _GEN_2636 : _GEN_2188; // @[Rob.scala 349:28]
  wire  _GEN_2845 = deq_ready_mask_0 ? _GEN_2637 : _GEN_2189; // @[Rob.scala 349:28]
  wire  _GEN_2846 = deq_ready_mask_0 ? _GEN_2638 : _GEN_2190; // @[Rob.scala 349:28]
  wire  _GEN_2847 = deq_ready_mask_0 ? _GEN_2639 : _GEN_2191; // @[Rob.scala 349:28]
  wire [5:0] _GEN_2848 = deq_ready_mask_0 ? _GEN_2640 : _GEN_1488; // @[Rob.scala 349:28]
  wire [5:0] _GEN_2849 = deq_ready_mask_0 ? _GEN_2641 : _GEN_1489; // @[Rob.scala 349:28]
  wire [5:0] _GEN_2850 = deq_ready_mask_0 ? _GEN_2642 : _GEN_1490; // @[Rob.scala 349:28]
  wire [5:0] _GEN_2851 = deq_ready_mask_0 ? _GEN_2643 : _GEN_1491; // @[Rob.scala 349:28]
  wire [5:0] _GEN_2852 = deq_ready_mask_0 ? _GEN_2644 : _GEN_1492; // @[Rob.scala 349:28]
  wire [5:0] _GEN_2853 = deq_ready_mask_0 ? _GEN_2645 : _GEN_1493; // @[Rob.scala 349:28]
  wire [5:0] _GEN_2854 = deq_ready_mask_0 ? _GEN_2646 : _GEN_1494; // @[Rob.scala 349:28]
  wire [5:0] _GEN_2855 = deq_ready_mask_0 ? _GEN_2647 : _GEN_1495; // @[Rob.scala 349:28]
  wire [2:0] _GEN_2856 = deq_ready_mask_0 ? _GEN_2648 : _GEN_1496; // @[Rob.scala 349:28]
  wire [2:0] _GEN_2857 = deq_ready_mask_0 ? _GEN_2649 : _GEN_1497; // @[Rob.scala 349:28]
  wire [2:0] _GEN_2858 = deq_ready_mask_0 ? _GEN_2650 : _GEN_1498; // @[Rob.scala 349:28]
  wire [2:0] _GEN_2859 = deq_ready_mask_0 ? _GEN_2651 : _GEN_1499; // @[Rob.scala 349:28]
  wire [2:0] _GEN_2860 = deq_ready_mask_0 ? _GEN_2652 : _GEN_1500; // @[Rob.scala 349:28]
  wire [2:0] _GEN_2861 = deq_ready_mask_0 ? _GEN_2653 : _GEN_1501; // @[Rob.scala 349:28]
  wire [2:0] _GEN_2862 = deq_ready_mask_0 ? _GEN_2654 : _GEN_1502; // @[Rob.scala 349:28]
  wire [2:0] _GEN_2863 = deq_ready_mask_0 ? _GEN_2655 : _GEN_1503; // @[Rob.scala 349:28]
  wire  _GEN_2864 = deq_ready_mask_0 ? _GEN_2656 : _GEN_1504; // @[Rob.scala 349:28]
  wire  _GEN_2865 = deq_ready_mask_0 ? _GEN_2657 : _GEN_1505; // @[Rob.scala 349:28]
  wire  _GEN_2866 = deq_ready_mask_0 ? _GEN_2658 : _GEN_1506; // @[Rob.scala 349:28]
  wire  _GEN_2867 = deq_ready_mask_0 ? _GEN_2659 : _GEN_1507; // @[Rob.scala 349:28]
  wire  _GEN_2868 = deq_ready_mask_0 ? _GEN_2660 : _GEN_1508; // @[Rob.scala 349:28]
  wire  _GEN_2869 = deq_ready_mask_0 ? _GEN_2661 : _GEN_1509; // @[Rob.scala 349:28]
  wire  _GEN_2870 = deq_ready_mask_0 ? _GEN_2662 : _GEN_1510; // @[Rob.scala 349:28]
  wire  _GEN_2871 = deq_ready_mask_0 ? _GEN_2663 : _GEN_1511; // @[Rob.scala 349:28]
  wire [31:0] _GEN_2872 = deq_ready_mask_0 ? _GEN_2664 : _GEN_1432; // @[Rob.scala 349:28]
  wire [31:0] _GEN_2873 = deq_ready_mask_0 ? _GEN_2665 : _GEN_1433; // @[Rob.scala 349:28]
  wire [31:0] _GEN_2874 = deq_ready_mask_0 ? _GEN_2666 : _GEN_1434; // @[Rob.scala 349:28]
  wire [31:0] _GEN_2875 = deq_ready_mask_0 ? _GEN_2667 : _GEN_1435; // @[Rob.scala 349:28]
  wire [31:0] _GEN_2876 = deq_ready_mask_0 ? _GEN_2668 : _GEN_1436; // @[Rob.scala 349:28]
  wire [31:0] _GEN_2877 = deq_ready_mask_0 ? _GEN_2669 : _GEN_1437; // @[Rob.scala 349:28]
  wire [31:0] _GEN_2878 = deq_ready_mask_0 ? _GEN_2670 : _GEN_1438; // @[Rob.scala 349:28]
  wire [31:0] _GEN_2879 = deq_ready_mask_0 ? _GEN_2671 : _GEN_1439; // @[Rob.scala 349:28]
  wire [4:0] _GEN_2880 = deq_ready_mask_0 ? _GEN_2672 : _GEN_1440; // @[Rob.scala 349:28]
  wire [4:0] _GEN_2881 = deq_ready_mask_0 ? _GEN_2673 : _GEN_1441; // @[Rob.scala 349:28]
  wire [4:0] _GEN_2882 = deq_ready_mask_0 ? _GEN_2674 : _GEN_1442; // @[Rob.scala 349:28]
  wire [4:0] _GEN_2883 = deq_ready_mask_0 ? _GEN_2675 : _GEN_1443; // @[Rob.scala 349:28]
  wire [4:0] _GEN_2884 = deq_ready_mask_0 ? _GEN_2676 : _GEN_1444; // @[Rob.scala 349:28]
  wire [4:0] _GEN_2885 = deq_ready_mask_0 ? _GEN_2677 : _GEN_1445; // @[Rob.scala 349:28]
  wire [4:0] _GEN_2886 = deq_ready_mask_0 ? _GEN_2678 : _GEN_1446; // @[Rob.scala 349:28]
  wire [4:0] _GEN_2887 = deq_ready_mask_0 ? _GEN_2679 : _GEN_1447; // @[Rob.scala 349:28]
  wire [31:0] _GEN_2888 = deq_ready_mask_0 ? _GEN_2680 : _GEN_2168; // @[Rob.scala 349:28]
  wire [31:0] _GEN_2889 = deq_ready_mask_0 ? _GEN_2681 : _GEN_2169; // @[Rob.scala 349:28]
  wire [31:0] _GEN_2890 = deq_ready_mask_0 ? _GEN_2682 : _GEN_2170; // @[Rob.scala 349:28]
  wire [31:0] _GEN_2891 = deq_ready_mask_0 ? _GEN_2683 : _GEN_2171; // @[Rob.scala 349:28]
  wire [31:0] _GEN_2892 = deq_ready_mask_0 ? _GEN_2684 : _GEN_2172; // @[Rob.scala 349:28]
  wire [31:0] _GEN_2893 = deq_ready_mask_0 ? _GEN_2685 : _GEN_2173; // @[Rob.scala 349:28]
  wire [31:0] _GEN_2894 = deq_ready_mask_0 ? _GEN_2686 : _GEN_2174; // @[Rob.scala 349:28]
  wire [31:0] _GEN_2895 = deq_ready_mask_0 ? _GEN_2687 : _GEN_2175; // @[Rob.scala 349:28]
  wire  _GEN_2904 = deq_ready_mask_0 ? _GEN_2696 : _GEN_2176; // @[Rob.scala 349:28]
  wire  _GEN_2905 = deq_ready_mask_0 ? _GEN_2697 : _GEN_2177; // @[Rob.scala 349:28]
  wire  _GEN_2906 = deq_ready_mask_0 ? _GEN_2698 : _GEN_2178; // @[Rob.scala 349:28]
  wire  _GEN_2907 = deq_ready_mask_0 ? _GEN_2699 : _GEN_2179; // @[Rob.scala 349:28]
  wire  _GEN_2908 = deq_ready_mask_0 ? _GEN_2700 : _GEN_2180; // @[Rob.scala 349:28]
  wire  _GEN_2909 = deq_ready_mask_0 ? _GEN_2701 : _GEN_2181; // @[Rob.scala 349:28]
  wire  _GEN_2910 = deq_ready_mask_0 ? _GEN_2702 : _GEN_2182; // @[Rob.scala 349:28]
  wire  _GEN_2911 = deq_ready_mask_0 ? _GEN_2703 : _GEN_2183; // @[Rob.scala 349:28]
  wire  _GEN_2920 = deq_ready_mask_0 ? _GEN_2712 : _GEN_1464; // @[Rob.scala 349:28]
  wire  _GEN_2921 = deq_ready_mask_0 ? _GEN_2713 : _GEN_1465; // @[Rob.scala 349:28]
  wire  _GEN_2922 = deq_ready_mask_0 ? _GEN_2714 : _GEN_1466; // @[Rob.scala 349:28]
  wire  _GEN_2923 = deq_ready_mask_0 ? _GEN_2715 : _GEN_1467; // @[Rob.scala 349:28]
  wire  _GEN_2924 = deq_ready_mask_0 ? _GEN_2716 : _GEN_1468; // @[Rob.scala 349:28]
  wire  _GEN_2925 = deq_ready_mask_0 ? _GEN_2717 : _GEN_1469; // @[Rob.scala 349:28]
  wire  _GEN_2926 = deq_ready_mask_0 ? _GEN_2718 : _GEN_1470; // @[Rob.scala 349:28]
  wire  _GEN_2927 = deq_ready_mask_0 ? _GEN_2719 : _GEN_1471; // @[Rob.scala 349:28]
  wire  _GEN_2936 = deq_ready_mask_0 ? _GEN_2728 : _GEN_1528; // @[Rob.scala 349:28]
  wire  _GEN_2937 = deq_ready_mask_0 ? _GEN_2729 : _GEN_1529; // @[Rob.scala 349:28]
  wire  _GEN_2938 = deq_ready_mask_0 ? _GEN_2730 : _GEN_1530; // @[Rob.scala 349:28]
  wire  _GEN_2939 = deq_ready_mask_0 ? _GEN_2731 : _GEN_1531; // @[Rob.scala 349:28]
  wire  _GEN_2940 = deq_ready_mask_0 ? _GEN_2732 : _GEN_1532; // @[Rob.scala 349:28]
  wire  _GEN_2941 = deq_ready_mask_0 ? _GEN_2733 : _GEN_1533; // @[Rob.scala 349:28]
  wire  _GEN_2942 = deq_ready_mask_0 ? _GEN_2734 : _GEN_1534; // @[Rob.scala 349:28]
  wire  _GEN_2943 = deq_ready_mask_0 ? _GEN_2735 : _GEN_1535; // @[Rob.scala 349:28]
  wire  _GEN_2944 = deq_ready_mask_0 ? _GEN_2736 : _GEN_2192; // @[Rob.scala 349:28]
  wire  _GEN_2945 = deq_ready_mask_0 ? _GEN_2737 : _GEN_2193; // @[Rob.scala 349:28]
  wire  _GEN_2946 = deq_ready_mask_0 ? _GEN_2738 : _GEN_2194; // @[Rob.scala 349:28]
  wire  _GEN_2947 = deq_ready_mask_0 ? _GEN_2739 : _GEN_2195; // @[Rob.scala 349:28]
  wire  _GEN_2948 = deq_ready_mask_0 ? _GEN_2740 : _GEN_2196; // @[Rob.scala 349:28]
  wire  _GEN_2949 = deq_ready_mask_0 ? _GEN_2741 : _GEN_2197; // @[Rob.scala 349:28]
  wire  _GEN_2950 = deq_ready_mask_0 ? _GEN_2742 : _GEN_2198; // @[Rob.scala 349:28]
  wire  _GEN_2951 = deq_ready_mask_0 ? _GEN_2743 : _GEN_2199; // @[Rob.scala 349:28]
  wire  _GEN_2952 = deq_ready_mask_0 ? _GEN_2744 : _GEN_2200; // @[Rob.scala 349:28]
  wire  _GEN_2953 = deq_ready_mask_0 ? _GEN_2745 : _GEN_2201; // @[Rob.scala 349:28]
  wire  _GEN_2954 = deq_ready_mask_0 ? _GEN_2746 : _GEN_2202; // @[Rob.scala 349:28]
  wire  _GEN_2955 = deq_ready_mask_0 ? _GEN_2747 : _GEN_2203; // @[Rob.scala 349:28]
  wire  _GEN_2956 = deq_ready_mask_0 ? _GEN_2748 : _GEN_2204; // @[Rob.scala 349:28]
  wire  _GEN_2957 = deq_ready_mask_0 ? _GEN_2749 : _GEN_2205; // @[Rob.scala 349:28]
  wire  _GEN_2958 = deq_ready_mask_0 ? _GEN_2750 : _GEN_2206; // @[Rob.scala 349:28]
  wire  _GEN_2959 = deq_ready_mask_0 ? _GEN_2751 : _GEN_2207; // @[Rob.scala 349:28]
  wire [3:0] _GEN_2960 = deq_ready_mask_0 ? _GEN_2752 : _GEN_1480; // @[Rob.scala 349:28]
  wire [3:0] _GEN_2961 = deq_ready_mask_0 ? _GEN_2753 : _GEN_1481; // @[Rob.scala 349:28]
  wire [3:0] _GEN_2962 = deq_ready_mask_0 ? _GEN_2754 : _GEN_1482; // @[Rob.scala 349:28]
  wire [3:0] _GEN_2963 = deq_ready_mask_0 ? _GEN_2755 : _GEN_1483; // @[Rob.scala 349:28]
  wire [3:0] _GEN_2964 = deq_ready_mask_0 ? _GEN_2756 : _GEN_1484; // @[Rob.scala 349:28]
  wire [3:0] _GEN_2965 = deq_ready_mask_0 ? _GEN_2757 : _GEN_1485; // @[Rob.scala 349:28]
  wire [3:0] _GEN_2966 = deq_ready_mask_0 ? _GEN_2758 : _GEN_1486; // @[Rob.scala 349:28]
  wire [3:0] _GEN_2967 = deq_ready_mask_0 ? _GEN_2759 : _GEN_1487; // @[Rob.scala 349:28]
  wire  _GEN_2968 = deq_ready_mask_0 ? _GEN_2760 : _GEN_2512; // @[Rob.scala 349:28]
  wire  _GEN_2969 = deq_ready_mask_0 ? _GEN_2761 : _GEN_2513; // @[Rob.scala 349:28]
  wire  _GEN_2970 = deq_ready_mask_0 ? _GEN_2762 : _GEN_2514; // @[Rob.scala 349:28]
  wire  _GEN_2971 = deq_ready_mask_0 ? _GEN_2763 : _GEN_2515; // @[Rob.scala 349:28]
  wire  _GEN_2972 = deq_ready_mask_0 ? _GEN_2764 : _GEN_2516; // @[Rob.scala 349:28]
  wire  _GEN_2973 = deq_ready_mask_0 ? _GEN_2765 : _GEN_2517; // @[Rob.scala 349:28]
  wire  _GEN_2974 = deq_ready_mask_0 ? _GEN_2766 : _GEN_2518; // @[Rob.scala 349:28]
  wire  _GEN_2975 = deq_ready_mask_0 ? _GEN_2767 : _GEN_2519; // @[Rob.scala 349:28]
  wire [2:0] _GEN_2976 = deq_ready_mask_0 ? _GEN_2768 : _GEN_2496; // @[Rob.scala 349:28]
  wire [2:0] _GEN_2977 = deq_ready_mask_0 ? _GEN_2769 : _GEN_2497; // @[Rob.scala 349:28]
  wire [2:0] _GEN_2978 = deq_ready_mask_0 ? _GEN_2770 : _GEN_2498; // @[Rob.scala 349:28]
  wire [2:0] _GEN_2979 = deq_ready_mask_0 ? _GEN_2771 : _GEN_2499; // @[Rob.scala 349:28]
  wire [2:0] _GEN_2980 = deq_ready_mask_0 ? _GEN_2772 : _GEN_2500; // @[Rob.scala 349:28]
  wire [2:0] _GEN_2981 = deq_ready_mask_0 ? _GEN_2773 : _GEN_2501; // @[Rob.scala 349:28]
  wire [2:0] _GEN_2982 = deq_ready_mask_0 ? _GEN_2774 : _GEN_2502; // @[Rob.scala 349:28]
  wire [2:0] _GEN_2983 = deq_ready_mask_0 ? _GEN_2775 : _GEN_2503; // @[Rob.scala 349:28]
  wire [31:0] _GEN_2984 = deq_ready_mask_0 ? _GEN_2776 : _GEN_2480; // @[Rob.scala 349:28]
  wire [31:0] _GEN_2985 = deq_ready_mask_0 ? _GEN_2777 : _GEN_2481; // @[Rob.scala 349:28]
  wire [31:0] _GEN_2986 = deq_ready_mask_0 ? _GEN_2778 : _GEN_2482; // @[Rob.scala 349:28]
  wire [31:0] _GEN_2987 = deq_ready_mask_0 ? _GEN_2779 : _GEN_2483; // @[Rob.scala 349:28]
  wire [31:0] _GEN_2988 = deq_ready_mask_0 ? _GEN_2780 : _GEN_2484; // @[Rob.scala 349:28]
  wire [31:0] _GEN_2989 = deq_ready_mask_0 ? _GEN_2781 : _GEN_2485; // @[Rob.scala 349:28]
  wire [31:0] _GEN_2990 = deq_ready_mask_0 ? _GEN_2782 : _GEN_2486; // @[Rob.scala 349:28]
  wire [31:0] _GEN_2991 = deq_ready_mask_0 ? _GEN_2783 : _GEN_2487; // @[Rob.scala 349:28]
  wire  _GEN_2992 = deq_ready_mask_0 ? _GEN_2784 : _GEN_2520; // @[Rob.scala 349:28]
  wire  _GEN_2993 = deq_ready_mask_0 ? _GEN_2785 : _GEN_2521; // @[Rob.scala 349:28]
  wire  _GEN_2994 = deq_ready_mask_0 ? _GEN_2786 : _GEN_2522; // @[Rob.scala 349:28]
  wire  _GEN_2995 = deq_ready_mask_0 ? _GEN_2787 : _GEN_2523; // @[Rob.scala 349:28]
  wire  _GEN_2996 = deq_ready_mask_0 ? _GEN_2788 : _GEN_2524; // @[Rob.scala 349:28]
  wire  _GEN_2997 = deq_ready_mask_0 ? _GEN_2789 : _GEN_2525; // @[Rob.scala 349:28]
  wire  _GEN_2998 = deq_ready_mask_0 ? _GEN_2790 : _GEN_2526; // @[Rob.scala 349:28]
  wire  _GEN_2999 = deq_ready_mask_0 ? _GEN_2791 : _GEN_2527; // @[Rob.scala 349:28]
  wire [2:0] _GEN_3000 = deq_ready_mask_0 ? _GEN_2792 : _GEN_2504; // @[Rob.scala 349:28]
  wire [2:0] _GEN_3001 = deq_ready_mask_0 ? _GEN_2793 : _GEN_2505; // @[Rob.scala 349:28]
  wire [2:0] _GEN_3002 = deq_ready_mask_0 ? _GEN_2794 : _GEN_2506; // @[Rob.scala 349:28]
  wire [2:0] _GEN_3003 = deq_ready_mask_0 ? _GEN_2795 : _GEN_2507; // @[Rob.scala 349:28]
  wire [2:0] _GEN_3004 = deq_ready_mask_0 ? _GEN_2796 : _GEN_2508; // @[Rob.scala 349:28]
  wire [2:0] _GEN_3005 = deq_ready_mask_0 ? _GEN_2797 : _GEN_2509; // @[Rob.scala 349:28]
  wire [2:0] _GEN_3006 = deq_ready_mask_0 ? _GEN_2798 : _GEN_2510; // @[Rob.scala 349:28]
  wire [2:0] _GEN_3007 = deq_ready_mask_0 ? _GEN_2799 : _GEN_2511; // @[Rob.scala 349:28]
  wire [31:0] _GEN_3008 = deq_ready_mask_0 ? _GEN_2800 : _GEN_2488; // @[Rob.scala 349:28]
  wire [31:0] _GEN_3009 = deq_ready_mask_0 ? _GEN_2801 : _GEN_2489; // @[Rob.scala 349:28]
  wire [31:0] _GEN_3010 = deq_ready_mask_0 ? _GEN_2802 : _GEN_2490; // @[Rob.scala 349:28]
  wire [31:0] _GEN_3011 = deq_ready_mask_0 ? _GEN_2803 : _GEN_2491; // @[Rob.scala 349:28]
  wire [31:0] _GEN_3012 = deq_ready_mask_0 ? _GEN_2804 : _GEN_2492; // @[Rob.scala 349:28]
  wire [31:0] _GEN_3013 = deq_ready_mask_0 ? _GEN_2805 : _GEN_2493; // @[Rob.scala 349:28]
  wire [31:0] _GEN_3014 = deq_ready_mask_0 ? _GEN_2806 : _GEN_2494; // @[Rob.scala 349:28]
  wire [31:0] _GEN_3015 = deq_ready_mask_0 ? _GEN_2807 : _GEN_2495; // @[Rob.scala 349:28]
  wire [31:0] _GEN_3016 = deq_ready_mask_0 ? _GEN_2808 : _GEN_2208; // @[Rob.scala 349:28]
  wire [31:0] _GEN_3017 = deq_ready_mask_0 ? _GEN_2809 : _GEN_2209; // @[Rob.scala 349:28]
  wire [31:0] _GEN_3018 = deq_ready_mask_0 ? _GEN_2810 : _GEN_2210; // @[Rob.scala 349:28]
  wire [31:0] _GEN_3019 = deq_ready_mask_0 ? _GEN_2811 : _GEN_2211; // @[Rob.scala 349:28]
  wire [31:0] _GEN_3020 = deq_ready_mask_0 ? _GEN_2812 : _GEN_2212; // @[Rob.scala 349:28]
  wire [31:0] _GEN_3021 = deq_ready_mask_0 ? _GEN_2813 : _GEN_2213; // @[Rob.scala 349:28]
  wire [31:0] _GEN_3022 = deq_ready_mask_0 ? _GEN_2814 : _GEN_2214; // @[Rob.scala 349:28]
  wire [31:0] _GEN_3023 = deq_ready_mask_0 ? _GEN_2815 : _GEN_2215; // @[Rob.scala 349:28]
  wire  _GEN_3024 = deq_ready_mask_0 ? _GEN_2816 : _GEN_2528; // @[Rob.scala 349:28]
  wire  _GEN_3025 = deq_ready_mask_0 ? _GEN_2817 : _GEN_2529; // @[Rob.scala 349:28]
  wire  _GEN_3026 = deq_ready_mask_0 ? _GEN_2818 : _GEN_2530; // @[Rob.scala 349:28]
  wire  _GEN_3027 = deq_ready_mask_0 ? _GEN_2819 : _GEN_2531; // @[Rob.scala 349:28]
  wire  _GEN_3028 = deq_ready_mask_0 ? _GEN_2820 : _GEN_2532; // @[Rob.scala 349:28]
  wire  _GEN_3029 = deq_ready_mask_0 ? _GEN_2821 : _GEN_2533; // @[Rob.scala 349:28]
  wire  _GEN_3030 = deq_ready_mask_0 ? _GEN_2822 : _GEN_2534; // @[Rob.scala 349:28]
  wire  _GEN_3031 = deq_ready_mask_0 ? _GEN_2823 : _GEN_2535; // @[Rob.scala 349:28]
  wire  _GEN_3032 = deq_ready_mask_0 ? _GEN_2824 : _GEN_1520; // @[Rob.scala 349:28]
  wire  _GEN_3033 = deq_ready_mask_0 ? _GEN_2825 : _GEN_1521; // @[Rob.scala 349:28]
  wire  _GEN_3034 = deq_ready_mask_0 ? _GEN_2826 : _GEN_1522; // @[Rob.scala 349:28]
  wire  _GEN_3035 = deq_ready_mask_0 ? _GEN_2827 : _GEN_1523; // @[Rob.scala 349:28]
  wire  _GEN_3036 = deq_ready_mask_0 ? _GEN_2828 : _GEN_1524; // @[Rob.scala 349:28]
  wire  _GEN_3037 = deq_ready_mask_0 ? _GEN_2829 : _GEN_1525; // @[Rob.scala 349:28]
  wire  _GEN_3038 = deq_ready_mask_0 ? _GEN_2830 : _GEN_1526; // @[Rob.scala 349:28]
  wire  _GEN_3039 = deq_ready_mask_0 ? _GEN_2831 : _GEN_1527; // @[Rob.scala 349:28]
  wire [31:0] _GEN_3041 = 3'h1 == dispatch_idxs_1 ? rob_info_1_commit_data : rob_info_0_commit_data; // @[Rob.scala 346:31 Rob.scala 346:31]
  wire [31:0] _GEN_3042 = 3'h2 == dispatch_idxs_1 ? rob_info_2_commit_data : _GEN_3041; // @[Rob.scala 346:31 Rob.scala 346:31]
  wire [31:0] _GEN_3043 = 3'h3 == dispatch_idxs_1 ? rob_info_3_commit_data : _GEN_3042; // @[Rob.scala 346:31 Rob.scala 346:31]
  wire [31:0] _GEN_3044 = 3'h4 == dispatch_idxs_1 ? rob_info_4_commit_data : _GEN_3043; // @[Rob.scala 346:31 Rob.scala 346:31]
  wire [31:0] _GEN_3045 = 3'h5 == dispatch_idxs_1 ? rob_info_5_commit_data : _GEN_3044; // @[Rob.scala 346:31 Rob.scala 346:31]
  wire [4:0] _GEN_3049 = 3'h1 == dispatch_idxs_1 ? rob_info_1_commit_addr : rob_info_0_commit_addr; // @[Rob.scala 348:31 Rob.scala 348:31]
  wire [4:0] _GEN_3050 = 3'h2 == dispatch_idxs_1 ? rob_info_2_commit_addr : _GEN_3049; // @[Rob.scala 348:31 Rob.scala 348:31]
  wire [4:0] _GEN_3051 = 3'h3 == dispatch_idxs_1 ? rob_info_3_commit_addr : _GEN_3050; // @[Rob.scala 348:31 Rob.scala 348:31]
  wire [4:0] _GEN_3052 = 3'h4 == dispatch_idxs_1 ? rob_info_4_commit_addr : _GEN_3051; // @[Rob.scala 348:31 Rob.scala 348:31]
  wire [4:0] _GEN_3053 = 3'h5 == dispatch_idxs_1 ? rob_info_5_commit_addr : _GEN_3052; // @[Rob.scala 348:31 Rob.scala 348:31]
  reg [31:0] branch_info_target_addr; // @[Rob.scala 385:24]
  reg [31:0] branch_info_inst_addr; // @[Rob.scala 385:24]
  reg [3:0] branch_info_gh_update; // @[Rob.scala 385:24]
  reg  branch_info_is_branch; // @[Rob.scala 385:24]
  reg  branch_info_is_taken; // @[Rob.scala 385:24]
  reg  branch_info_predict_miss; // @[Rob.scala 385:24]
  reg  branch_info_valid; // @[Rob.scala 386:34]
  wire [2:0] _GEN_3529 = flush_idx ? dispatch_idxs_1 : dispatch_idxs_0; // @[Rob.scala 388:27 Rob.scala 388:27]
  wire [31:0] _GEN_3531 = 3'h1 == _GEN_3529 ? rob_info_1_imm_data : rob_info_0_imm_data; // @[Rob.scala 388:27 Rob.scala 388:27]
  wire [31:0] _GEN_3532 = 3'h2 == _GEN_3529 ? rob_info_2_imm_data : _GEN_3531; // @[Rob.scala 388:27 Rob.scala 388:27]
  wire [31:0] _GEN_3533 = 3'h3 == _GEN_3529 ? rob_info_3_imm_data : _GEN_3532; // @[Rob.scala 388:27 Rob.scala 388:27]
  wire [31:0] _GEN_3534 = 3'h4 == _GEN_3529 ? rob_info_4_imm_data : _GEN_3533; // @[Rob.scala 388:27 Rob.scala 388:27]
  wire [31:0] _GEN_3535 = 3'h5 == _GEN_3529 ? rob_info_5_imm_data : _GEN_3534; // @[Rob.scala 388:27 Rob.scala 388:27]
  wire [31:0] _GEN_3536 = 3'h6 == _GEN_3529 ? rob_info_6_imm_data : _GEN_3535; // @[Rob.scala 388:27 Rob.scala 388:27]
  wire [31:0] _GEN_3539 = 3'h1 == _GEN_3529 ? rob_info_1_inst_addr : rob_info_0_inst_addr; // @[Rob.scala 389:25 Rob.scala 389:25]
  wire [31:0] _GEN_3540 = 3'h2 == _GEN_3529 ? rob_info_2_inst_addr : _GEN_3539; // @[Rob.scala 389:25 Rob.scala 389:25]
  wire [31:0] _GEN_3541 = 3'h3 == _GEN_3529 ? rob_info_3_inst_addr : _GEN_3540; // @[Rob.scala 389:25 Rob.scala 389:25]
  wire [31:0] _GEN_3542 = 3'h4 == _GEN_3529 ? rob_info_4_inst_addr : _GEN_3541; // @[Rob.scala 389:25 Rob.scala 389:25]
  wire [31:0] _GEN_3543 = 3'h5 == _GEN_3529 ? rob_info_5_inst_addr : _GEN_3542; // @[Rob.scala 389:25 Rob.scala 389:25]
  wire [31:0] _GEN_3544 = 3'h6 == _GEN_3529 ? rob_info_6_inst_addr : _GEN_3543; // @[Rob.scala 389:25 Rob.scala 389:25]
  wire [3:0] _GEN_3547 = 3'h1 == _GEN_3529 ? rob_info_1_gh_info : rob_info_0_gh_info; // @[Rob.scala 390:25 Rob.scala 390:25]
  wire [3:0] _GEN_3548 = 3'h2 == _GEN_3529 ? rob_info_2_gh_info : _GEN_3547; // @[Rob.scala 390:25 Rob.scala 390:25]
  wire [3:0] _GEN_3549 = 3'h3 == _GEN_3529 ? rob_info_3_gh_info : _GEN_3548; // @[Rob.scala 390:25 Rob.scala 390:25]
  wire [3:0] _GEN_3550 = 3'h4 == _GEN_3529 ? rob_info_4_gh_info : _GEN_3549; // @[Rob.scala 390:25 Rob.scala 390:25]
  wire [3:0] _GEN_3551 = 3'h5 == _GEN_3529 ? rob_info_5_gh_info : _GEN_3550; // @[Rob.scala 390:25 Rob.scala 390:25]
  wire [3:0] _GEN_3552 = 3'h6 == _GEN_3529 ? rob_info_6_gh_info : _GEN_3551; // @[Rob.scala 390:25 Rob.scala 390:25]
  wire  _GEN_3555 = 3'h1 == _GEN_3529 ? rob_info_1_is_branch : rob_info_0_is_branch; // @[Rob.scala 391:25 Rob.scala 391:25]
  wire  _GEN_3556 = 3'h2 == _GEN_3529 ? rob_info_2_is_branch : _GEN_3555; // @[Rob.scala 391:25 Rob.scala 391:25]
  wire  _GEN_3557 = 3'h3 == _GEN_3529 ? rob_info_3_is_branch : _GEN_3556; // @[Rob.scala 391:25 Rob.scala 391:25]
  wire  _GEN_3558 = 3'h4 == _GEN_3529 ? rob_info_4_is_branch : _GEN_3557; // @[Rob.scala 391:25 Rob.scala 391:25]
  wire  _GEN_3559 = 3'h5 == _GEN_3529 ? rob_info_5_is_branch : _GEN_3558; // @[Rob.scala 391:25 Rob.scala 391:25]
  wire  _GEN_3560 = 3'h6 == _GEN_3529 ? rob_info_6_is_branch : _GEN_3559; // @[Rob.scala 391:25 Rob.scala 391:25]
  wire  _GEN_3563 = 3'h1 == _GEN_3529 ? rob_info_1_is_taken : rob_info_0_is_taken; // @[Rob.scala 392:24 Rob.scala 392:24]
  wire  _GEN_3564 = 3'h2 == _GEN_3529 ? rob_info_2_is_taken : _GEN_3563; // @[Rob.scala 392:24 Rob.scala 392:24]
  wire  _GEN_3565 = 3'h3 == _GEN_3529 ? rob_info_3_is_taken : _GEN_3564; // @[Rob.scala 392:24 Rob.scala 392:24]
  wire  _GEN_3566 = 3'h4 == _GEN_3529 ? rob_info_4_is_taken : _GEN_3565; // @[Rob.scala 392:24 Rob.scala 392:24]
  wire  _GEN_3567 = 3'h5 == _GEN_3529 ? rob_info_5_is_taken : _GEN_3566; // @[Rob.scala 392:24 Rob.scala 392:24]
  wire  _GEN_3568 = 3'h6 == _GEN_3529 ? rob_info_6_is_taken : _GEN_3567; // @[Rob.scala 392:24 Rob.scala 392:24]
  wire  _GEN_3571 = 3'h1 == _GEN_3529 ? rob_info_1_predict_miss : rob_info_0_predict_miss; // @[Rob.scala 393:28 Rob.scala 393:28]
  wire  _GEN_3572 = 3'h2 == _GEN_3529 ? rob_info_2_predict_miss : _GEN_3571; // @[Rob.scala 393:28 Rob.scala 393:28]
  wire  _GEN_3573 = 3'h3 == _GEN_3529 ? rob_info_3_predict_miss : _GEN_3572; // @[Rob.scala 393:28 Rob.scala 393:28]
  wire  _GEN_3574 = 3'h4 == _GEN_3529 ? rob_info_4_predict_miss : _GEN_3573; // @[Rob.scala 393:28 Rob.scala 393:28]
  wire  _GEN_3575 = 3'h5 == _GEN_3529 ? rob_info_5_predict_miss : _GEN_3574; // @[Rob.scala 393:28 Rob.scala 393:28]
  wire  _GEN_3576 = 3'h6 == _GEN_3529 ? rob_info_6_predict_miss : _GEN_3575; // @[Rob.scala 393:28 Rob.scala 393:28]
  wire  _GEN_3578 = deq_ready_mask_0 ? 1'h0 : maybe_full; // @[Rob.scala 402:22 Rob.scala 403:16 Rob.scala 179:31]
  wire  _GEN_3579 = do_enq | _GEN_3578; // @[Rob.scala 400:16 Rob.scala 401:16]
  wire  _GEN_3580 = flush | waiting_delay; // @[Rob.scala 411:15 Rob.scala 412:19 Rob.scala 187:30]
  wire  _GEN_3591 = waiting_delay & deq_ready_mask_0; // @[Rob.scala 429:22 Rob.scala 440:15]
  assign io_rob_allocate_allocate_resp_valid = enq_valid_mask_0 | enq_valid_mask_1; // @[Rob.scala 198:43]
  assign io_rob_allocate_allocate_resp_bits_rob_idx_0 = {hi_3,lo_5}; // @[Cat.scala 30:58]
  assign io_rob_allocate_allocate_resp_bits_rob_idx_1 = {hi_7,lo_9}; // @[Cat.scala 30:58]
  assign io_rob_allocate_allocate_resp_bits_enq_valid_mask_0 = _T_4 & inst_valid_mask_0; // @[Rob.scala 197:79]
  assign io_rob_allocate_allocate_resp_bits_enq_valid_mask_1 = _T_11 & inst_valid_mask_1; // @[Rob.scala 197:79]
  assign io_dispatch_info_o_0_valid = _GEN_391 & _GEN_399; // @[Rob.scala 224:50]
  assign io_dispatch_info_o_0_bits_uop = 3'h7 == _GEN_407 ? rob_info_7_uop : _GEN_414; // @[Rob.scala 227:36 Rob.scala 227:36]
  assign io_dispatch_info_o_0_bits_need_imm = 3'h7 == _GEN_407 ? rob_info_7_need_imm : _GEN_422; // @[Rob.scala 228:41 Rob.scala 228:41]
  assign io_dispatch_info_o_0_bits_rob_idx = 3'h7 == dispatch_idx ? dispatch_idxs_7 : _GEN_406; // @[Rob.scala 226:40 Rob.scala 226:40]
  assign io_dispatch_info_o_0_bits_op1_data = 3'h7 == _GEN_407 ? rob_info_7_op1_data : _GEN_438; // @[Rob.scala 230:41 Rob.scala 230:41]
  assign io_dispatch_info_o_0_bits_op2_data = 3'h7 == _GEN_407 ? rob_info_7_op2_data : _GEN_446; // @[Rob.scala 231:41 Rob.scala 231:41]
  assign io_dispatch_info_o_0_bits_imm_data = 3'h7 == _GEN_407 ? rob_info_7_imm_data : _GEN_454; // @[Rob.scala 232:41 Rob.scala 232:41]
  assign io_dispatch_info_o_1_valid = _GEN_487 & _GEN_495; // @[Rob.scala 224:50]
  assign io_dispatch_info_o_1_bits_uop = 3'h7 == _GEN_503 ? rob_info_7_uop : _GEN_510; // @[Rob.scala 227:36 Rob.scala 227:36]
  assign io_dispatch_info_o_1_bits_need_imm = 3'h7 == _GEN_503 ? rob_info_7_need_imm : _GEN_518; // @[Rob.scala 228:41 Rob.scala 228:41]
  assign io_dispatch_info_o_1_bits_rob_idx = 3'h7 == dispatch_idx_1 ? dispatch_idxs_7 : _GEN_502; // @[Rob.scala 226:40 Rob.scala 226:40]
  assign io_dispatch_info_o_1_bits_op1_data = 3'h7 == _GEN_503 ? rob_info_7_op1_data : _GEN_534; // @[Rob.scala 230:41 Rob.scala 230:41]
  assign io_dispatch_info_o_1_bits_op2_data = 3'h7 == _GEN_503 ? rob_info_7_op2_data : _GEN_542; // @[Rob.scala 231:41 Rob.scala 231:41]
  assign io_dispatch_info_o_1_bits_imm_data = 3'h7 == _GEN_503 ? rob_info_7_imm_data : _GEN_550; // @[Rob.scala 232:41 Rob.scala 232:41]
  assign io_dispatch_info_o_2_valid = _GEN_583 & _GEN_591; // @[Rob.scala 224:50]
  assign io_dispatch_info_o_2_bits_uop = 3'h7 == _GEN_599 ? rob_info_7_uop : _GEN_606; // @[Rob.scala 227:36 Rob.scala 227:36]
  assign io_dispatch_info_o_2_bits_rob_idx = 3'h7 == dispatch_idx_2 ? dispatch_idxs_7 : _GEN_598; // @[Rob.scala 226:40 Rob.scala 226:40]
  assign io_dispatch_info_o_2_bits_inst_addr = 3'h7 == _GEN_599 ? rob_info_7_inst_addr : _GEN_622; // @[Rob.scala 229:42 Rob.scala 229:42]
  assign io_dispatch_info_o_2_bits_op1_data = 3'h7 == _GEN_599 ? rob_info_7_op1_data : _GEN_630; // @[Rob.scala 230:41 Rob.scala 230:41]
  assign io_dispatch_info_o_2_bits_op2_data = 3'h7 == _GEN_599 ? rob_info_7_op2_data : _GEN_638; // @[Rob.scala 231:41 Rob.scala 231:41]
  assign io_dispatch_info_o_2_bits_imm_data = 3'h7 == _GEN_599 ? rob_info_7_imm_data : _GEN_646; // @[Rob.scala 232:41 Rob.scala 232:41]
  assign io_dispatch_info_o_2_bits_predict_taken = 3'h7 == _GEN_599 ? rob_info_7_predict_taken : _GEN_654; // @[Rob.scala 233:46 Rob.scala 233:46]
  assign io_dispatch_info_o_3_valid = _GEN_679 & _GEN_687; // @[Rob.scala 224:50]
  assign io_dispatch_info_o_3_bits_rob_idx = 3'h7 == dispatch_idx_3 ? dispatch_idxs_7 : _GEN_694; // @[Rob.scala 226:40 Rob.scala 226:40]
  assign io_dispatch_info_o_3_bits_op1_data = 3'h7 == _GEN_695 ? rob_info_7_op1_data : _GEN_726; // @[Rob.scala 230:41 Rob.scala 230:41]
  assign io_dispatch_info_o_3_bits_op2_data = 3'h7 == _GEN_695 ? rob_info_7_op2_data : _GEN_734; // @[Rob.scala 231:41 Rob.scala 231:41]
  assign io_dispatch_info_o_4_valid = _GEN_775 & _GEN_783; // @[Rob.scala 224:50]
  assign io_dispatch_info_o_4_bits_uop = 3'h7 == _GEN_791 ? rob_info_7_uop : _GEN_798; // @[Rob.scala 227:36 Rob.scala 227:36]
  assign io_dispatch_info_o_4_bits_rob_idx = 3'h7 == dispatch_idx_4 ? dispatch_idxs_7 : _GEN_790; // @[Rob.scala 226:40 Rob.scala 226:40]
  assign io_dispatch_info_o_4_bits_op1_data = 3'h7 == _GEN_791 ? rob_info_7_op1_data : _GEN_822; // @[Rob.scala 230:41 Rob.scala 230:41]
  assign io_dispatch_info_o_4_bits_op2_data = 3'h7 == _GEN_791 ? rob_info_7_op2_data : _GEN_830; // @[Rob.scala 231:41 Rob.scala 231:41]
  assign io_dispatch_info_o_4_bits_imm_data = 3'h7 == _GEN_791 ? rob_info_7_imm_data : _GEN_838; // @[Rob.scala 232:41 Rob.scala 232:41]
  assign io_rob_commit_0_valid = rob_commit_valid_0; // @[Rob.scala 353:27]
  assign io_rob_commit_0_bits_des_rob = rob_commit_0_des_rob; // @[Rob.scala 352:26]
  assign io_rob_commit_0_bits_commit_addr = rob_commit_0_commit_addr; // @[Rob.scala 352:26]
  assign io_rob_commit_0_bits_commit_data = rob_commit_0_commit_data; // @[Rob.scala 352:26]
  assign io_rob_commit_1_valid = rob_commit_valid_1; // @[Rob.scala 353:27]
  assign io_rob_commit_1_bits_des_rob = rob_commit_1_des_rob; // @[Rob.scala 352:26]
  assign io_rob_commit_1_bits_commit_addr = rob_commit_1_commit_addr; // @[Rob.scala 352:26]
  assign io_rob_commit_1_bits_commit_data = rob_commit_1_commit_data; // @[Rob.scala 352:26]
  assign io_branch_info_valid = branch_info_valid; // @[Rob.scala 396:23]
  assign io_branch_info_bits_target_addr = branch_info_target_addr; // @[Rob.scala 395:22]
  assign io_branch_info_bits_inst_addr = branch_info_inst_addr; // @[Rob.scala 395:22]
  assign io_branch_info_bits_gh_update = branch_info_gh_update; // @[Rob.scala 395:22]
  assign io_branch_info_bits_is_branch = branch_info_is_branch; // @[Rob.scala 395:22]
  assign io_branch_info_bits_is_taken = branch_info_is_taken; // @[Rob.scala 395:22]
  assign io_branch_info_bits_predict_miss = branch_info_predict_miss; // @[Rob.scala 395:22]
  assign io_need_flush = need_flush; // @[Rob.scala 443:16]
  always @(posedge clock) begin
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_0_is_valid <= 1'h0; // @[Rob.scala 42:13]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_0_is_valid <= 1'h0; // @[Rob.scala 42:13]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h0 == dispatch_idxs_1) begin // @[Rob.scala 42:13]
        rob_info_0_is_valid <= 1'h0; // @[Rob.scala 42:13]
      end else begin
        rob_info_0_is_valid <= _GEN_2832;
      end
    end else begin
      rob_info_0_is_valid <= _GEN_2832;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_0_busy <= 1'h0; // @[Rob.scala 43:9]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_0_busy <= 1'h0; // @[Rob.scala 43:9]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h0 == dispatch_idxs_1) begin // @[Rob.scala 43:9]
        rob_info_0_busy <= 1'h0; // @[Rob.scala 43:9]
      end else begin
        rob_info_0_busy <= _GEN_2840;
      end
    end else begin
      rob_info_0_busy <= _GEN_2840;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_0_uop <= 6'h0; // @[Rob.scala 44:8]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_0_uop <= 6'h0; // @[Rob.scala 44:8]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h0 == dispatch_idxs_1) begin // @[Rob.scala 44:8]
        rob_info_0_uop <= 6'h0; // @[Rob.scala 44:8]
      end else begin
        rob_info_0_uop <= _GEN_2848;
      end
    end else begin
      rob_info_0_uop <= _GEN_2848;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_0_unit_sel <= 3'h0; // @[Rob.scala 45:13]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_0_unit_sel <= 3'h0; // @[Rob.scala 45:13]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h0 == dispatch_idxs_1) begin // @[Rob.scala 45:13]
        rob_info_0_unit_sel <= 3'h0; // @[Rob.scala 45:13]
      end else begin
        rob_info_0_unit_sel <= _GEN_2856;
      end
    end else begin
      rob_info_0_unit_sel <= _GEN_2856;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_0_need_imm <= 1'h0; // @[Rob.scala 46:13]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_0_need_imm <= 1'h0; // @[Rob.scala 46:13]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h0 == dispatch_idxs_1) begin // @[Rob.scala 46:13]
        rob_info_0_need_imm <= 1'h0; // @[Rob.scala 46:13]
      end else begin
        rob_info_0_need_imm <= _GEN_2864;
      end
    end else begin
      rob_info_0_need_imm <= _GEN_2864;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_0_inst_addr <= 32'h0; // @[Rob.scala 47:14]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_0_inst_addr <= 32'h0; // @[Rob.scala 47:14]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h0 == dispatch_idxs_1) begin // @[Rob.scala 47:14]
        rob_info_0_inst_addr <= 32'h0; // @[Rob.scala 47:14]
      end else begin
        rob_info_0_inst_addr <= _GEN_2872;
      end
    end else begin
      rob_info_0_inst_addr <= _GEN_2872;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_0_commit_addr <= 5'h0; // @[Rob.scala 48:16]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_0_commit_addr <= 5'h0; // @[Rob.scala 48:16]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h0 == dispatch_idxs_1) begin // @[Rob.scala 48:16]
        rob_info_0_commit_addr <= 5'h0; // @[Rob.scala 48:16]
      end else begin
        rob_info_0_commit_addr <= _GEN_2880;
      end
    end else begin
      rob_info_0_commit_addr <= _GEN_2880;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_0_commit_data <= 32'h0; // @[Rob.scala 49:16]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_0_commit_data <= 32'h0; // @[Rob.scala 49:16]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h0 == dispatch_idxs_1) begin // @[Rob.scala 49:16]
        rob_info_0_commit_data <= 32'h0; // @[Rob.scala 49:16]
      end else begin
        rob_info_0_commit_data <= _GEN_2888;
      end
    end else begin
      rob_info_0_commit_data <= _GEN_2888;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_0_commit_ready <= 1'h0; // @[Rob.scala 51:17]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_0_commit_ready <= 1'h0; // @[Rob.scala 51:17]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h0 == dispatch_idxs_1) begin // @[Rob.scala 51:17]
        rob_info_0_commit_ready <= 1'h0; // @[Rob.scala 51:17]
      end else begin
        rob_info_0_commit_ready <= _GEN_2904;
      end
    end else begin
      rob_info_0_commit_ready <= _GEN_2904;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_0_is_branch <= 1'h0; // @[Rob.scala 53:14]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_0_is_branch <= 1'h0; // @[Rob.scala 53:14]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h0 == dispatch_idxs_1) begin // @[Rob.scala 53:14]
        rob_info_0_is_branch <= 1'h0; // @[Rob.scala 53:14]
      end else begin
        rob_info_0_is_branch <= _GEN_2920;
      end
    end else begin
      rob_info_0_is_branch <= _GEN_2920;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_0_predict_taken <= 1'h0; // @[Rob.scala 55:18]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_0_predict_taken <= 1'h0; // @[Rob.scala 55:18]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h0 == dispatch_idxs_1) begin // @[Rob.scala 55:18]
        rob_info_0_predict_taken <= 1'h0; // @[Rob.scala 55:18]
      end else begin
        rob_info_0_predict_taken <= _GEN_2936;
      end
    end else begin
      rob_info_0_predict_taken <= _GEN_2936;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_0_is_taken <= 1'h0; // @[Rob.scala 56:13]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_0_is_taken <= 1'h0; // @[Rob.scala 56:13]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h0 == dispatch_idxs_1) begin // @[Rob.scala 56:13]
        rob_info_0_is_taken <= 1'h0; // @[Rob.scala 56:13]
      end else begin
        rob_info_0_is_taken <= _GEN_2944;
      end
    end else begin
      rob_info_0_is_taken <= _GEN_2944;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_0_predict_miss <= 1'h0; // @[Rob.scala 57:17]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_0_predict_miss <= 1'h0; // @[Rob.scala 57:17]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h0 == dispatch_idxs_1) begin // @[Rob.scala 57:17]
        rob_info_0_predict_miss <= 1'h0; // @[Rob.scala 57:17]
      end else begin
        rob_info_0_predict_miss <= _GEN_2952;
      end
    end else begin
      rob_info_0_predict_miss <= _GEN_2952;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_0_gh_info <= 4'h0; // @[Rob.scala 58:12]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_0_gh_info <= 4'h0; // @[Rob.scala 58:12]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h0 == dispatch_idxs_1) begin // @[Rob.scala 58:12]
        rob_info_0_gh_info <= 4'h0; // @[Rob.scala 58:12]
      end else begin
        rob_info_0_gh_info <= _GEN_2960;
      end
    end else begin
      rob_info_0_gh_info <= _GEN_2960;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_0_op1_ready <= 1'h0; // @[Rob.scala 59:14]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_0_op1_ready <= 1'h0; // @[Rob.scala 59:14]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h0 == dispatch_idxs_1) begin // @[Rob.scala 59:14]
        rob_info_0_op1_ready <= 1'h0; // @[Rob.scala 59:14]
      end else begin
        rob_info_0_op1_ready <= _GEN_2968;
      end
    end else begin
      rob_info_0_op1_ready <= _GEN_2968;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_0_op1_tag <= 3'h0; // @[Rob.scala 60:12]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_0_op1_tag <= 3'h0; // @[Rob.scala 60:12]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h0 == dispatch_idxs_1) begin // @[Rob.scala 60:12]
        rob_info_0_op1_tag <= 3'h0; // @[Rob.scala 60:12]
      end else begin
        rob_info_0_op1_tag <= _GEN_2976;
      end
    end else begin
      rob_info_0_op1_tag <= _GEN_2976;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_0_op1_data <= 32'h0; // @[Rob.scala 61:13]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_0_op1_data <= 32'h0; // @[Rob.scala 61:13]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h0 == dispatch_idxs_1) begin // @[Rob.scala 61:13]
        rob_info_0_op1_data <= 32'h0; // @[Rob.scala 61:13]
      end else begin
        rob_info_0_op1_data <= _GEN_2984;
      end
    end else begin
      rob_info_0_op1_data <= _GEN_2984;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_0_op2_ready <= 1'h0; // @[Rob.scala 62:14]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_0_op2_ready <= 1'h0; // @[Rob.scala 62:14]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h0 == dispatch_idxs_1) begin // @[Rob.scala 62:14]
        rob_info_0_op2_ready <= 1'h0; // @[Rob.scala 62:14]
      end else begin
        rob_info_0_op2_ready <= _GEN_2992;
      end
    end else begin
      rob_info_0_op2_ready <= _GEN_2992;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_0_op2_tag <= 3'h0; // @[Rob.scala 63:12]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_0_op2_tag <= 3'h0; // @[Rob.scala 63:12]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h0 == dispatch_idxs_1) begin // @[Rob.scala 63:12]
        rob_info_0_op2_tag <= 3'h0; // @[Rob.scala 63:12]
      end else begin
        rob_info_0_op2_tag <= _GEN_3000;
      end
    end else begin
      rob_info_0_op2_tag <= _GEN_3000;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_0_op2_data <= 32'h0; // @[Rob.scala 64:13]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_0_op2_data <= 32'h0; // @[Rob.scala 64:13]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h0 == dispatch_idxs_1) begin // @[Rob.scala 64:13]
        rob_info_0_op2_data <= 32'h0; // @[Rob.scala 64:13]
      end else begin
        rob_info_0_op2_data <= _GEN_3008;
      end
    end else begin
      rob_info_0_op2_data <= _GEN_3008;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_0_imm_data <= 32'h0; // @[Rob.scala 65:13]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_0_imm_data <= 32'h0; // @[Rob.scala 65:13]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h0 == dispatch_idxs_1) begin // @[Rob.scala 65:13]
        rob_info_0_imm_data <= 32'h0; // @[Rob.scala 65:13]
      end else begin
        rob_info_0_imm_data <= _GEN_3016;
      end
    end else begin
      rob_info_0_imm_data <= _GEN_3016;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_0_is_init <= 1'h0; // @[Rob.scala 66:13]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_0_is_init <= 1'h0; // @[Rob.scala 66:13]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h0 == dispatch_idxs_1) begin // @[Rob.scala 66:13]
        rob_info_0_is_init <= 1'h0; // @[Rob.scala 66:13]
      end else begin
        rob_info_0_is_init <= _GEN_3024;
      end
    end else begin
      rob_info_0_is_init <= _GEN_3024;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_0_flush_on_commit <= 1'h0; // @[Rob.scala 67:20]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_0_flush_on_commit <= 1'h0; // @[Rob.scala 67:20]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h0 == dispatch_idxs_1) begin // @[Rob.scala 67:20]
        rob_info_0_flush_on_commit <= 1'h0; // @[Rob.scala 67:20]
      end else begin
        rob_info_0_flush_on_commit <= _GEN_3032;
      end
    end else begin
      rob_info_0_flush_on_commit <= _GEN_3032;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_1_is_valid <= 1'h0; // @[Rob.scala 42:13]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_1_is_valid <= 1'h0; // @[Rob.scala 42:13]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h1 == dispatch_idxs_1) begin // @[Rob.scala 42:13]
        rob_info_1_is_valid <= 1'h0; // @[Rob.scala 42:13]
      end else begin
        rob_info_1_is_valid <= _GEN_2833;
      end
    end else begin
      rob_info_1_is_valid <= _GEN_2833;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_1_busy <= 1'h0; // @[Rob.scala 43:9]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_1_busy <= 1'h0; // @[Rob.scala 43:9]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h1 == dispatch_idxs_1) begin // @[Rob.scala 43:9]
        rob_info_1_busy <= 1'h0; // @[Rob.scala 43:9]
      end else begin
        rob_info_1_busy <= _GEN_2841;
      end
    end else begin
      rob_info_1_busy <= _GEN_2841;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_1_uop <= 6'h0; // @[Rob.scala 44:8]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_1_uop <= 6'h0; // @[Rob.scala 44:8]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h1 == dispatch_idxs_1) begin // @[Rob.scala 44:8]
        rob_info_1_uop <= 6'h0; // @[Rob.scala 44:8]
      end else begin
        rob_info_1_uop <= _GEN_2849;
      end
    end else begin
      rob_info_1_uop <= _GEN_2849;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_1_unit_sel <= 3'h0; // @[Rob.scala 45:13]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_1_unit_sel <= 3'h0; // @[Rob.scala 45:13]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h1 == dispatch_idxs_1) begin // @[Rob.scala 45:13]
        rob_info_1_unit_sel <= 3'h0; // @[Rob.scala 45:13]
      end else begin
        rob_info_1_unit_sel <= _GEN_2857;
      end
    end else begin
      rob_info_1_unit_sel <= _GEN_2857;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_1_need_imm <= 1'h0; // @[Rob.scala 46:13]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_1_need_imm <= 1'h0; // @[Rob.scala 46:13]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h1 == dispatch_idxs_1) begin // @[Rob.scala 46:13]
        rob_info_1_need_imm <= 1'h0; // @[Rob.scala 46:13]
      end else begin
        rob_info_1_need_imm <= _GEN_2865;
      end
    end else begin
      rob_info_1_need_imm <= _GEN_2865;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_1_inst_addr <= 32'h0; // @[Rob.scala 47:14]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_1_inst_addr <= 32'h0; // @[Rob.scala 47:14]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h1 == dispatch_idxs_1) begin // @[Rob.scala 47:14]
        rob_info_1_inst_addr <= 32'h0; // @[Rob.scala 47:14]
      end else begin
        rob_info_1_inst_addr <= _GEN_2873;
      end
    end else begin
      rob_info_1_inst_addr <= _GEN_2873;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_1_commit_addr <= 5'h0; // @[Rob.scala 48:16]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_1_commit_addr <= 5'h0; // @[Rob.scala 48:16]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h1 == dispatch_idxs_1) begin // @[Rob.scala 48:16]
        rob_info_1_commit_addr <= 5'h0; // @[Rob.scala 48:16]
      end else begin
        rob_info_1_commit_addr <= _GEN_2881;
      end
    end else begin
      rob_info_1_commit_addr <= _GEN_2881;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_1_commit_data <= 32'h0; // @[Rob.scala 49:16]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_1_commit_data <= 32'h0; // @[Rob.scala 49:16]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h1 == dispatch_idxs_1) begin // @[Rob.scala 49:16]
        rob_info_1_commit_data <= 32'h0; // @[Rob.scala 49:16]
      end else begin
        rob_info_1_commit_data <= _GEN_2889;
      end
    end else begin
      rob_info_1_commit_data <= _GEN_2889;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_1_commit_ready <= 1'h0; // @[Rob.scala 51:17]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_1_commit_ready <= 1'h0; // @[Rob.scala 51:17]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h1 == dispatch_idxs_1) begin // @[Rob.scala 51:17]
        rob_info_1_commit_ready <= 1'h0; // @[Rob.scala 51:17]
      end else begin
        rob_info_1_commit_ready <= _GEN_2905;
      end
    end else begin
      rob_info_1_commit_ready <= _GEN_2905;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_1_is_branch <= 1'h0; // @[Rob.scala 53:14]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_1_is_branch <= 1'h0; // @[Rob.scala 53:14]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h1 == dispatch_idxs_1) begin // @[Rob.scala 53:14]
        rob_info_1_is_branch <= 1'h0; // @[Rob.scala 53:14]
      end else begin
        rob_info_1_is_branch <= _GEN_2921;
      end
    end else begin
      rob_info_1_is_branch <= _GEN_2921;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_1_predict_taken <= 1'h0; // @[Rob.scala 55:18]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_1_predict_taken <= 1'h0; // @[Rob.scala 55:18]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h1 == dispatch_idxs_1) begin // @[Rob.scala 55:18]
        rob_info_1_predict_taken <= 1'h0; // @[Rob.scala 55:18]
      end else begin
        rob_info_1_predict_taken <= _GEN_2937;
      end
    end else begin
      rob_info_1_predict_taken <= _GEN_2937;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_1_is_taken <= 1'h0; // @[Rob.scala 56:13]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_1_is_taken <= 1'h0; // @[Rob.scala 56:13]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h1 == dispatch_idxs_1) begin // @[Rob.scala 56:13]
        rob_info_1_is_taken <= 1'h0; // @[Rob.scala 56:13]
      end else begin
        rob_info_1_is_taken <= _GEN_2945;
      end
    end else begin
      rob_info_1_is_taken <= _GEN_2945;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_1_predict_miss <= 1'h0; // @[Rob.scala 57:17]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_1_predict_miss <= 1'h0; // @[Rob.scala 57:17]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h1 == dispatch_idxs_1) begin // @[Rob.scala 57:17]
        rob_info_1_predict_miss <= 1'h0; // @[Rob.scala 57:17]
      end else begin
        rob_info_1_predict_miss <= _GEN_2953;
      end
    end else begin
      rob_info_1_predict_miss <= _GEN_2953;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_1_gh_info <= 4'h0; // @[Rob.scala 58:12]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_1_gh_info <= 4'h0; // @[Rob.scala 58:12]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h1 == dispatch_idxs_1) begin // @[Rob.scala 58:12]
        rob_info_1_gh_info <= 4'h0; // @[Rob.scala 58:12]
      end else begin
        rob_info_1_gh_info <= _GEN_2961;
      end
    end else begin
      rob_info_1_gh_info <= _GEN_2961;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_1_op1_ready <= 1'h0; // @[Rob.scala 59:14]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_1_op1_ready <= 1'h0; // @[Rob.scala 59:14]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h1 == dispatch_idxs_1) begin // @[Rob.scala 59:14]
        rob_info_1_op1_ready <= 1'h0; // @[Rob.scala 59:14]
      end else begin
        rob_info_1_op1_ready <= _GEN_2969;
      end
    end else begin
      rob_info_1_op1_ready <= _GEN_2969;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_1_op1_tag <= 3'h0; // @[Rob.scala 60:12]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_1_op1_tag <= 3'h0; // @[Rob.scala 60:12]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h1 == dispatch_idxs_1) begin // @[Rob.scala 60:12]
        rob_info_1_op1_tag <= 3'h0; // @[Rob.scala 60:12]
      end else begin
        rob_info_1_op1_tag <= _GEN_2977;
      end
    end else begin
      rob_info_1_op1_tag <= _GEN_2977;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_1_op1_data <= 32'h0; // @[Rob.scala 61:13]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_1_op1_data <= 32'h0; // @[Rob.scala 61:13]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h1 == dispatch_idxs_1) begin // @[Rob.scala 61:13]
        rob_info_1_op1_data <= 32'h0; // @[Rob.scala 61:13]
      end else begin
        rob_info_1_op1_data <= _GEN_2985;
      end
    end else begin
      rob_info_1_op1_data <= _GEN_2985;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_1_op2_ready <= 1'h0; // @[Rob.scala 62:14]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_1_op2_ready <= 1'h0; // @[Rob.scala 62:14]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h1 == dispatch_idxs_1) begin // @[Rob.scala 62:14]
        rob_info_1_op2_ready <= 1'h0; // @[Rob.scala 62:14]
      end else begin
        rob_info_1_op2_ready <= _GEN_2993;
      end
    end else begin
      rob_info_1_op2_ready <= _GEN_2993;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_1_op2_tag <= 3'h0; // @[Rob.scala 63:12]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_1_op2_tag <= 3'h0; // @[Rob.scala 63:12]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h1 == dispatch_idxs_1) begin // @[Rob.scala 63:12]
        rob_info_1_op2_tag <= 3'h0; // @[Rob.scala 63:12]
      end else begin
        rob_info_1_op2_tag <= _GEN_3001;
      end
    end else begin
      rob_info_1_op2_tag <= _GEN_3001;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_1_op2_data <= 32'h0; // @[Rob.scala 64:13]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_1_op2_data <= 32'h0; // @[Rob.scala 64:13]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h1 == dispatch_idxs_1) begin // @[Rob.scala 64:13]
        rob_info_1_op2_data <= 32'h0; // @[Rob.scala 64:13]
      end else begin
        rob_info_1_op2_data <= _GEN_3009;
      end
    end else begin
      rob_info_1_op2_data <= _GEN_3009;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_1_imm_data <= 32'h0; // @[Rob.scala 65:13]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_1_imm_data <= 32'h0; // @[Rob.scala 65:13]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h1 == dispatch_idxs_1) begin // @[Rob.scala 65:13]
        rob_info_1_imm_data <= 32'h0; // @[Rob.scala 65:13]
      end else begin
        rob_info_1_imm_data <= _GEN_3017;
      end
    end else begin
      rob_info_1_imm_data <= _GEN_3017;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_1_is_init <= 1'h0; // @[Rob.scala 66:13]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_1_is_init <= 1'h0; // @[Rob.scala 66:13]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h1 == dispatch_idxs_1) begin // @[Rob.scala 66:13]
        rob_info_1_is_init <= 1'h0; // @[Rob.scala 66:13]
      end else begin
        rob_info_1_is_init <= _GEN_3025;
      end
    end else begin
      rob_info_1_is_init <= _GEN_3025;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_1_flush_on_commit <= 1'h0; // @[Rob.scala 67:20]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_1_flush_on_commit <= 1'h0; // @[Rob.scala 67:20]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h1 == dispatch_idxs_1) begin // @[Rob.scala 67:20]
        rob_info_1_flush_on_commit <= 1'h0; // @[Rob.scala 67:20]
      end else begin
        rob_info_1_flush_on_commit <= _GEN_3033;
      end
    end else begin
      rob_info_1_flush_on_commit <= _GEN_3033;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_2_is_valid <= 1'h0; // @[Rob.scala 42:13]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_2_is_valid <= 1'h0; // @[Rob.scala 42:13]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h2 == dispatch_idxs_1) begin // @[Rob.scala 42:13]
        rob_info_2_is_valid <= 1'h0; // @[Rob.scala 42:13]
      end else begin
        rob_info_2_is_valid <= _GEN_2834;
      end
    end else begin
      rob_info_2_is_valid <= _GEN_2834;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_2_busy <= 1'h0; // @[Rob.scala 43:9]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_2_busy <= 1'h0; // @[Rob.scala 43:9]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h2 == dispatch_idxs_1) begin // @[Rob.scala 43:9]
        rob_info_2_busy <= 1'h0; // @[Rob.scala 43:9]
      end else begin
        rob_info_2_busy <= _GEN_2842;
      end
    end else begin
      rob_info_2_busy <= _GEN_2842;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_2_uop <= 6'h0; // @[Rob.scala 44:8]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_2_uop <= 6'h0; // @[Rob.scala 44:8]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h2 == dispatch_idxs_1) begin // @[Rob.scala 44:8]
        rob_info_2_uop <= 6'h0; // @[Rob.scala 44:8]
      end else begin
        rob_info_2_uop <= _GEN_2850;
      end
    end else begin
      rob_info_2_uop <= _GEN_2850;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_2_unit_sel <= 3'h0; // @[Rob.scala 45:13]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_2_unit_sel <= 3'h0; // @[Rob.scala 45:13]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h2 == dispatch_idxs_1) begin // @[Rob.scala 45:13]
        rob_info_2_unit_sel <= 3'h0; // @[Rob.scala 45:13]
      end else begin
        rob_info_2_unit_sel <= _GEN_2858;
      end
    end else begin
      rob_info_2_unit_sel <= _GEN_2858;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_2_need_imm <= 1'h0; // @[Rob.scala 46:13]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_2_need_imm <= 1'h0; // @[Rob.scala 46:13]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h2 == dispatch_idxs_1) begin // @[Rob.scala 46:13]
        rob_info_2_need_imm <= 1'h0; // @[Rob.scala 46:13]
      end else begin
        rob_info_2_need_imm <= _GEN_2866;
      end
    end else begin
      rob_info_2_need_imm <= _GEN_2866;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_2_inst_addr <= 32'h0; // @[Rob.scala 47:14]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_2_inst_addr <= 32'h0; // @[Rob.scala 47:14]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h2 == dispatch_idxs_1) begin // @[Rob.scala 47:14]
        rob_info_2_inst_addr <= 32'h0; // @[Rob.scala 47:14]
      end else begin
        rob_info_2_inst_addr <= _GEN_2874;
      end
    end else begin
      rob_info_2_inst_addr <= _GEN_2874;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_2_commit_addr <= 5'h0; // @[Rob.scala 48:16]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_2_commit_addr <= 5'h0; // @[Rob.scala 48:16]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h2 == dispatch_idxs_1) begin // @[Rob.scala 48:16]
        rob_info_2_commit_addr <= 5'h0; // @[Rob.scala 48:16]
      end else begin
        rob_info_2_commit_addr <= _GEN_2882;
      end
    end else begin
      rob_info_2_commit_addr <= _GEN_2882;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_2_commit_data <= 32'h0; // @[Rob.scala 49:16]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_2_commit_data <= 32'h0; // @[Rob.scala 49:16]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h2 == dispatch_idxs_1) begin // @[Rob.scala 49:16]
        rob_info_2_commit_data <= 32'h0; // @[Rob.scala 49:16]
      end else begin
        rob_info_2_commit_data <= _GEN_2890;
      end
    end else begin
      rob_info_2_commit_data <= _GEN_2890;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_2_commit_ready <= 1'h0; // @[Rob.scala 51:17]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_2_commit_ready <= 1'h0; // @[Rob.scala 51:17]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h2 == dispatch_idxs_1) begin // @[Rob.scala 51:17]
        rob_info_2_commit_ready <= 1'h0; // @[Rob.scala 51:17]
      end else begin
        rob_info_2_commit_ready <= _GEN_2906;
      end
    end else begin
      rob_info_2_commit_ready <= _GEN_2906;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_2_is_branch <= 1'h0; // @[Rob.scala 53:14]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_2_is_branch <= 1'h0; // @[Rob.scala 53:14]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h2 == dispatch_idxs_1) begin // @[Rob.scala 53:14]
        rob_info_2_is_branch <= 1'h0; // @[Rob.scala 53:14]
      end else begin
        rob_info_2_is_branch <= _GEN_2922;
      end
    end else begin
      rob_info_2_is_branch <= _GEN_2922;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_2_predict_taken <= 1'h0; // @[Rob.scala 55:18]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_2_predict_taken <= 1'h0; // @[Rob.scala 55:18]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h2 == dispatch_idxs_1) begin // @[Rob.scala 55:18]
        rob_info_2_predict_taken <= 1'h0; // @[Rob.scala 55:18]
      end else begin
        rob_info_2_predict_taken <= _GEN_2938;
      end
    end else begin
      rob_info_2_predict_taken <= _GEN_2938;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_2_is_taken <= 1'h0; // @[Rob.scala 56:13]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_2_is_taken <= 1'h0; // @[Rob.scala 56:13]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h2 == dispatch_idxs_1) begin // @[Rob.scala 56:13]
        rob_info_2_is_taken <= 1'h0; // @[Rob.scala 56:13]
      end else begin
        rob_info_2_is_taken <= _GEN_2946;
      end
    end else begin
      rob_info_2_is_taken <= _GEN_2946;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_2_predict_miss <= 1'h0; // @[Rob.scala 57:17]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_2_predict_miss <= 1'h0; // @[Rob.scala 57:17]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h2 == dispatch_idxs_1) begin // @[Rob.scala 57:17]
        rob_info_2_predict_miss <= 1'h0; // @[Rob.scala 57:17]
      end else begin
        rob_info_2_predict_miss <= _GEN_2954;
      end
    end else begin
      rob_info_2_predict_miss <= _GEN_2954;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_2_gh_info <= 4'h0; // @[Rob.scala 58:12]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_2_gh_info <= 4'h0; // @[Rob.scala 58:12]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h2 == dispatch_idxs_1) begin // @[Rob.scala 58:12]
        rob_info_2_gh_info <= 4'h0; // @[Rob.scala 58:12]
      end else begin
        rob_info_2_gh_info <= _GEN_2962;
      end
    end else begin
      rob_info_2_gh_info <= _GEN_2962;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_2_op1_ready <= 1'h0; // @[Rob.scala 59:14]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_2_op1_ready <= 1'h0; // @[Rob.scala 59:14]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h2 == dispatch_idxs_1) begin // @[Rob.scala 59:14]
        rob_info_2_op1_ready <= 1'h0; // @[Rob.scala 59:14]
      end else begin
        rob_info_2_op1_ready <= _GEN_2970;
      end
    end else begin
      rob_info_2_op1_ready <= _GEN_2970;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_2_op1_tag <= 3'h0; // @[Rob.scala 60:12]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_2_op1_tag <= 3'h0; // @[Rob.scala 60:12]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h2 == dispatch_idxs_1) begin // @[Rob.scala 60:12]
        rob_info_2_op1_tag <= 3'h0; // @[Rob.scala 60:12]
      end else begin
        rob_info_2_op1_tag <= _GEN_2978;
      end
    end else begin
      rob_info_2_op1_tag <= _GEN_2978;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_2_op1_data <= 32'h0; // @[Rob.scala 61:13]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_2_op1_data <= 32'h0; // @[Rob.scala 61:13]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h2 == dispatch_idxs_1) begin // @[Rob.scala 61:13]
        rob_info_2_op1_data <= 32'h0; // @[Rob.scala 61:13]
      end else begin
        rob_info_2_op1_data <= _GEN_2986;
      end
    end else begin
      rob_info_2_op1_data <= _GEN_2986;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_2_op2_ready <= 1'h0; // @[Rob.scala 62:14]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_2_op2_ready <= 1'h0; // @[Rob.scala 62:14]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h2 == dispatch_idxs_1) begin // @[Rob.scala 62:14]
        rob_info_2_op2_ready <= 1'h0; // @[Rob.scala 62:14]
      end else begin
        rob_info_2_op2_ready <= _GEN_2994;
      end
    end else begin
      rob_info_2_op2_ready <= _GEN_2994;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_2_op2_tag <= 3'h0; // @[Rob.scala 63:12]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_2_op2_tag <= 3'h0; // @[Rob.scala 63:12]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h2 == dispatch_idxs_1) begin // @[Rob.scala 63:12]
        rob_info_2_op2_tag <= 3'h0; // @[Rob.scala 63:12]
      end else begin
        rob_info_2_op2_tag <= _GEN_3002;
      end
    end else begin
      rob_info_2_op2_tag <= _GEN_3002;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_2_op2_data <= 32'h0; // @[Rob.scala 64:13]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_2_op2_data <= 32'h0; // @[Rob.scala 64:13]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h2 == dispatch_idxs_1) begin // @[Rob.scala 64:13]
        rob_info_2_op2_data <= 32'h0; // @[Rob.scala 64:13]
      end else begin
        rob_info_2_op2_data <= _GEN_3010;
      end
    end else begin
      rob_info_2_op2_data <= _GEN_3010;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_2_imm_data <= 32'h0; // @[Rob.scala 65:13]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_2_imm_data <= 32'h0; // @[Rob.scala 65:13]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h2 == dispatch_idxs_1) begin // @[Rob.scala 65:13]
        rob_info_2_imm_data <= 32'h0; // @[Rob.scala 65:13]
      end else begin
        rob_info_2_imm_data <= _GEN_3018;
      end
    end else begin
      rob_info_2_imm_data <= _GEN_3018;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_2_is_init <= 1'h0; // @[Rob.scala 66:13]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_2_is_init <= 1'h0; // @[Rob.scala 66:13]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h2 == dispatch_idxs_1) begin // @[Rob.scala 66:13]
        rob_info_2_is_init <= 1'h0; // @[Rob.scala 66:13]
      end else begin
        rob_info_2_is_init <= _GEN_3026;
      end
    end else begin
      rob_info_2_is_init <= _GEN_3026;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_2_flush_on_commit <= 1'h0; // @[Rob.scala 67:20]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_2_flush_on_commit <= 1'h0; // @[Rob.scala 67:20]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h2 == dispatch_idxs_1) begin // @[Rob.scala 67:20]
        rob_info_2_flush_on_commit <= 1'h0; // @[Rob.scala 67:20]
      end else begin
        rob_info_2_flush_on_commit <= _GEN_3034;
      end
    end else begin
      rob_info_2_flush_on_commit <= _GEN_3034;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_3_is_valid <= 1'h0; // @[Rob.scala 42:13]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_3_is_valid <= 1'h0; // @[Rob.scala 42:13]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h3 == dispatch_idxs_1) begin // @[Rob.scala 42:13]
        rob_info_3_is_valid <= 1'h0; // @[Rob.scala 42:13]
      end else begin
        rob_info_3_is_valid <= _GEN_2835;
      end
    end else begin
      rob_info_3_is_valid <= _GEN_2835;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_3_busy <= 1'h0; // @[Rob.scala 43:9]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_3_busy <= 1'h0; // @[Rob.scala 43:9]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h3 == dispatch_idxs_1) begin // @[Rob.scala 43:9]
        rob_info_3_busy <= 1'h0; // @[Rob.scala 43:9]
      end else begin
        rob_info_3_busy <= _GEN_2843;
      end
    end else begin
      rob_info_3_busy <= _GEN_2843;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_3_uop <= 6'h0; // @[Rob.scala 44:8]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_3_uop <= 6'h0; // @[Rob.scala 44:8]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h3 == dispatch_idxs_1) begin // @[Rob.scala 44:8]
        rob_info_3_uop <= 6'h0; // @[Rob.scala 44:8]
      end else begin
        rob_info_3_uop <= _GEN_2851;
      end
    end else begin
      rob_info_3_uop <= _GEN_2851;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_3_unit_sel <= 3'h0; // @[Rob.scala 45:13]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_3_unit_sel <= 3'h0; // @[Rob.scala 45:13]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h3 == dispatch_idxs_1) begin // @[Rob.scala 45:13]
        rob_info_3_unit_sel <= 3'h0; // @[Rob.scala 45:13]
      end else begin
        rob_info_3_unit_sel <= _GEN_2859;
      end
    end else begin
      rob_info_3_unit_sel <= _GEN_2859;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_3_need_imm <= 1'h0; // @[Rob.scala 46:13]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_3_need_imm <= 1'h0; // @[Rob.scala 46:13]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h3 == dispatch_idxs_1) begin // @[Rob.scala 46:13]
        rob_info_3_need_imm <= 1'h0; // @[Rob.scala 46:13]
      end else begin
        rob_info_3_need_imm <= _GEN_2867;
      end
    end else begin
      rob_info_3_need_imm <= _GEN_2867;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_3_inst_addr <= 32'h0; // @[Rob.scala 47:14]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_3_inst_addr <= 32'h0; // @[Rob.scala 47:14]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h3 == dispatch_idxs_1) begin // @[Rob.scala 47:14]
        rob_info_3_inst_addr <= 32'h0; // @[Rob.scala 47:14]
      end else begin
        rob_info_3_inst_addr <= _GEN_2875;
      end
    end else begin
      rob_info_3_inst_addr <= _GEN_2875;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_3_commit_addr <= 5'h0; // @[Rob.scala 48:16]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_3_commit_addr <= 5'h0; // @[Rob.scala 48:16]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h3 == dispatch_idxs_1) begin // @[Rob.scala 48:16]
        rob_info_3_commit_addr <= 5'h0; // @[Rob.scala 48:16]
      end else begin
        rob_info_3_commit_addr <= _GEN_2883;
      end
    end else begin
      rob_info_3_commit_addr <= _GEN_2883;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_3_commit_data <= 32'h0; // @[Rob.scala 49:16]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_3_commit_data <= 32'h0; // @[Rob.scala 49:16]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h3 == dispatch_idxs_1) begin // @[Rob.scala 49:16]
        rob_info_3_commit_data <= 32'h0; // @[Rob.scala 49:16]
      end else begin
        rob_info_3_commit_data <= _GEN_2891;
      end
    end else begin
      rob_info_3_commit_data <= _GEN_2891;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_3_commit_ready <= 1'h0; // @[Rob.scala 51:17]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_3_commit_ready <= 1'h0; // @[Rob.scala 51:17]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h3 == dispatch_idxs_1) begin // @[Rob.scala 51:17]
        rob_info_3_commit_ready <= 1'h0; // @[Rob.scala 51:17]
      end else begin
        rob_info_3_commit_ready <= _GEN_2907;
      end
    end else begin
      rob_info_3_commit_ready <= _GEN_2907;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_3_is_branch <= 1'h0; // @[Rob.scala 53:14]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_3_is_branch <= 1'h0; // @[Rob.scala 53:14]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h3 == dispatch_idxs_1) begin // @[Rob.scala 53:14]
        rob_info_3_is_branch <= 1'h0; // @[Rob.scala 53:14]
      end else begin
        rob_info_3_is_branch <= _GEN_2923;
      end
    end else begin
      rob_info_3_is_branch <= _GEN_2923;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_3_predict_taken <= 1'h0; // @[Rob.scala 55:18]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_3_predict_taken <= 1'h0; // @[Rob.scala 55:18]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h3 == dispatch_idxs_1) begin // @[Rob.scala 55:18]
        rob_info_3_predict_taken <= 1'h0; // @[Rob.scala 55:18]
      end else begin
        rob_info_3_predict_taken <= _GEN_2939;
      end
    end else begin
      rob_info_3_predict_taken <= _GEN_2939;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_3_is_taken <= 1'h0; // @[Rob.scala 56:13]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_3_is_taken <= 1'h0; // @[Rob.scala 56:13]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h3 == dispatch_idxs_1) begin // @[Rob.scala 56:13]
        rob_info_3_is_taken <= 1'h0; // @[Rob.scala 56:13]
      end else begin
        rob_info_3_is_taken <= _GEN_2947;
      end
    end else begin
      rob_info_3_is_taken <= _GEN_2947;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_3_predict_miss <= 1'h0; // @[Rob.scala 57:17]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_3_predict_miss <= 1'h0; // @[Rob.scala 57:17]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h3 == dispatch_idxs_1) begin // @[Rob.scala 57:17]
        rob_info_3_predict_miss <= 1'h0; // @[Rob.scala 57:17]
      end else begin
        rob_info_3_predict_miss <= _GEN_2955;
      end
    end else begin
      rob_info_3_predict_miss <= _GEN_2955;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_3_gh_info <= 4'h0; // @[Rob.scala 58:12]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_3_gh_info <= 4'h0; // @[Rob.scala 58:12]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h3 == dispatch_idxs_1) begin // @[Rob.scala 58:12]
        rob_info_3_gh_info <= 4'h0; // @[Rob.scala 58:12]
      end else begin
        rob_info_3_gh_info <= _GEN_2963;
      end
    end else begin
      rob_info_3_gh_info <= _GEN_2963;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_3_op1_ready <= 1'h0; // @[Rob.scala 59:14]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_3_op1_ready <= 1'h0; // @[Rob.scala 59:14]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h3 == dispatch_idxs_1) begin // @[Rob.scala 59:14]
        rob_info_3_op1_ready <= 1'h0; // @[Rob.scala 59:14]
      end else begin
        rob_info_3_op1_ready <= _GEN_2971;
      end
    end else begin
      rob_info_3_op1_ready <= _GEN_2971;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_3_op1_tag <= 3'h0; // @[Rob.scala 60:12]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_3_op1_tag <= 3'h0; // @[Rob.scala 60:12]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h3 == dispatch_idxs_1) begin // @[Rob.scala 60:12]
        rob_info_3_op1_tag <= 3'h0; // @[Rob.scala 60:12]
      end else begin
        rob_info_3_op1_tag <= _GEN_2979;
      end
    end else begin
      rob_info_3_op1_tag <= _GEN_2979;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_3_op1_data <= 32'h0; // @[Rob.scala 61:13]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_3_op1_data <= 32'h0; // @[Rob.scala 61:13]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h3 == dispatch_idxs_1) begin // @[Rob.scala 61:13]
        rob_info_3_op1_data <= 32'h0; // @[Rob.scala 61:13]
      end else begin
        rob_info_3_op1_data <= _GEN_2987;
      end
    end else begin
      rob_info_3_op1_data <= _GEN_2987;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_3_op2_ready <= 1'h0; // @[Rob.scala 62:14]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_3_op2_ready <= 1'h0; // @[Rob.scala 62:14]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h3 == dispatch_idxs_1) begin // @[Rob.scala 62:14]
        rob_info_3_op2_ready <= 1'h0; // @[Rob.scala 62:14]
      end else begin
        rob_info_3_op2_ready <= _GEN_2995;
      end
    end else begin
      rob_info_3_op2_ready <= _GEN_2995;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_3_op2_tag <= 3'h0; // @[Rob.scala 63:12]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_3_op2_tag <= 3'h0; // @[Rob.scala 63:12]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h3 == dispatch_idxs_1) begin // @[Rob.scala 63:12]
        rob_info_3_op2_tag <= 3'h0; // @[Rob.scala 63:12]
      end else begin
        rob_info_3_op2_tag <= _GEN_3003;
      end
    end else begin
      rob_info_3_op2_tag <= _GEN_3003;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_3_op2_data <= 32'h0; // @[Rob.scala 64:13]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_3_op2_data <= 32'h0; // @[Rob.scala 64:13]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h3 == dispatch_idxs_1) begin // @[Rob.scala 64:13]
        rob_info_3_op2_data <= 32'h0; // @[Rob.scala 64:13]
      end else begin
        rob_info_3_op2_data <= _GEN_3011;
      end
    end else begin
      rob_info_3_op2_data <= _GEN_3011;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_3_imm_data <= 32'h0; // @[Rob.scala 65:13]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_3_imm_data <= 32'h0; // @[Rob.scala 65:13]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h3 == dispatch_idxs_1) begin // @[Rob.scala 65:13]
        rob_info_3_imm_data <= 32'h0; // @[Rob.scala 65:13]
      end else begin
        rob_info_3_imm_data <= _GEN_3019;
      end
    end else begin
      rob_info_3_imm_data <= _GEN_3019;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_3_is_init <= 1'h0; // @[Rob.scala 66:13]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_3_is_init <= 1'h0; // @[Rob.scala 66:13]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h3 == dispatch_idxs_1) begin // @[Rob.scala 66:13]
        rob_info_3_is_init <= 1'h0; // @[Rob.scala 66:13]
      end else begin
        rob_info_3_is_init <= _GEN_3027;
      end
    end else begin
      rob_info_3_is_init <= _GEN_3027;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_3_flush_on_commit <= 1'h0; // @[Rob.scala 67:20]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_3_flush_on_commit <= 1'h0; // @[Rob.scala 67:20]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h3 == dispatch_idxs_1) begin // @[Rob.scala 67:20]
        rob_info_3_flush_on_commit <= 1'h0; // @[Rob.scala 67:20]
      end else begin
        rob_info_3_flush_on_commit <= _GEN_3035;
      end
    end else begin
      rob_info_3_flush_on_commit <= _GEN_3035;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_4_is_valid <= 1'h0; // @[Rob.scala 42:13]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_4_is_valid <= 1'h0; // @[Rob.scala 42:13]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h4 == dispatch_idxs_1) begin // @[Rob.scala 42:13]
        rob_info_4_is_valid <= 1'h0; // @[Rob.scala 42:13]
      end else begin
        rob_info_4_is_valid <= _GEN_2836;
      end
    end else begin
      rob_info_4_is_valid <= _GEN_2836;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_4_busy <= 1'h0; // @[Rob.scala 43:9]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_4_busy <= 1'h0; // @[Rob.scala 43:9]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h4 == dispatch_idxs_1) begin // @[Rob.scala 43:9]
        rob_info_4_busy <= 1'h0; // @[Rob.scala 43:9]
      end else begin
        rob_info_4_busy <= _GEN_2844;
      end
    end else begin
      rob_info_4_busy <= _GEN_2844;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_4_uop <= 6'h0; // @[Rob.scala 44:8]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_4_uop <= 6'h0; // @[Rob.scala 44:8]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h4 == dispatch_idxs_1) begin // @[Rob.scala 44:8]
        rob_info_4_uop <= 6'h0; // @[Rob.scala 44:8]
      end else begin
        rob_info_4_uop <= _GEN_2852;
      end
    end else begin
      rob_info_4_uop <= _GEN_2852;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_4_unit_sel <= 3'h0; // @[Rob.scala 45:13]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_4_unit_sel <= 3'h0; // @[Rob.scala 45:13]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h4 == dispatch_idxs_1) begin // @[Rob.scala 45:13]
        rob_info_4_unit_sel <= 3'h0; // @[Rob.scala 45:13]
      end else begin
        rob_info_4_unit_sel <= _GEN_2860;
      end
    end else begin
      rob_info_4_unit_sel <= _GEN_2860;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_4_need_imm <= 1'h0; // @[Rob.scala 46:13]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_4_need_imm <= 1'h0; // @[Rob.scala 46:13]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h4 == dispatch_idxs_1) begin // @[Rob.scala 46:13]
        rob_info_4_need_imm <= 1'h0; // @[Rob.scala 46:13]
      end else begin
        rob_info_4_need_imm <= _GEN_2868;
      end
    end else begin
      rob_info_4_need_imm <= _GEN_2868;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_4_inst_addr <= 32'h0; // @[Rob.scala 47:14]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_4_inst_addr <= 32'h0; // @[Rob.scala 47:14]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h4 == dispatch_idxs_1) begin // @[Rob.scala 47:14]
        rob_info_4_inst_addr <= 32'h0; // @[Rob.scala 47:14]
      end else begin
        rob_info_4_inst_addr <= _GEN_2876;
      end
    end else begin
      rob_info_4_inst_addr <= _GEN_2876;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_4_commit_addr <= 5'h0; // @[Rob.scala 48:16]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_4_commit_addr <= 5'h0; // @[Rob.scala 48:16]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h4 == dispatch_idxs_1) begin // @[Rob.scala 48:16]
        rob_info_4_commit_addr <= 5'h0; // @[Rob.scala 48:16]
      end else begin
        rob_info_4_commit_addr <= _GEN_2884;
      end
    end else begin
      rob_info_4_commit_addr <= _GEN_2884;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_4_commit_data <= 32'h0; // @[Rob.scala 49:16]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_4_commit_data <= 32'h0; // @[Rob.scala 49:16]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h4 == dispatch_idxs_1) begin // @[Rob.scala 49:16]
        rob_info_4_commit_data <= 32'h0; // @[Rob.scala 49:16]
      end else begin
        rob_info_4_commit_data <= _GEN_2892;
      end
    end else begin
      rob_info_4_commit_data <= _GEN_2892;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_4_commit_ready <= 1'h0; // @[Rob.scala 51:17]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_4_commit_ready <= 1'h0; // @[Rob.scala 51:17]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h4 == dispatch_idxs_1) begin // @[Rob.scala 51:17]
        rob_info_4_commit_ready <= 1'h0; // @[Rob.scala 51:17]
      end else begin
        rob_info_4_commit_ready <= _GEN_2908;
      end
    end else begin
      rob_info_4_commit_ready <= _GEN_2908;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_4_is_branch <= 1'h0; // @[Rob.scala 53:14]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_4_is_branch <= 1'h0; // @[Rob.scala 53:14]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h4 == dispatch_idxs_1) begin // @[Rob.scala 53:14]
        rob_info_4_is_branch <= 1'h0; // @[Rob.scala 53:14]
      end else begin
        rob_info_4_is_branch <= _GEN_2924;
      end
    end else begin
      rob_info_4_is_branch <= _GEN_2924;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_4_predict_taken <= 1'h0; // @[Rob.scala 55:18]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_4_predict_taken <= 1'h0; // @[Rob.scala 55:18]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h4 == dispatch_idxs_1) begin // @[Rob.scala 55:18]
        rob_info_4_predict_taken <= 1'h0; // @[Rob.scala 55:18]
      end else begin
        rob_info_4_predict_taken <= _GEN_2940;
      end
    end else begin
      rob_info_4_predict_taken <= _GEN_2940;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_4_is_taken <= 1'h0; // @[Rob.scala 56:13]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_4_is_taken <= 1'h0; // @[Rob.scala 56:13]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h4 == dispatch_idxs_1) begin // @[Rob.scala 56:13]
        rob_info_4_is_taken <= 1'h0; // @[Rob.scala 56:13]
      end else begin
        rob_info_4_is_taken <= _GEN_2948;
      end
    end else begin
      rob_info_4_is_taken <= _GEN_2948;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_4_predict_miss <= 1'h0; // @[Rob.scala 57:17]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_4_predict_miss <= 1'h0; // @[Rob.scala 57:17]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h4 == dispatch_idxs_1) begin // @[Rob.scala 57:17]
        rob_info_4_predict_miss <= 1'h0; // @[Rob.scala 57:17]
      end else begin
        rob_info_4_predict_miss <= _GEN_2956;
      end
    end else begin
      rob_info_4_predict_miss <= _GEN_2956;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_4_gh_info <= 4'h0; // @[Rob.scala 58:12]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_4_gh_info <= 4'h0; // @[Rob.scala 58:12]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h4 == dispatch_idxs_1) begin // @[Rob.scala 58:12]
        rob_info_4_gh_info <= 4'h0; // @[Rob.scala 58:12]
      end else begin
        rob_info_4_gh_info <= _GEN_2964;
      end
    end else begin
      rob_info_4_gh_info <= _GEN_2964;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_4_op1_ready <= 1'h0; // @[Rob.scala 59:14]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_4_op1_ready <= 1'h0; // @[Rob.scala 59:14]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h4 == dispatch_idxs_1) begin // @[Rob.scala 59:14]
        rob_info_4_op1_ready <= 1'h0; // @[Rob.scala 59:14]
      end else begin
        rob_info_4_op1_ready <= _GEN_2972;
      end
    end else begin
      rob_info_4_op1_ready <= _GEN_2972;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_4_op1_tag <= 3'h0; // @[Rob.scala 60:12]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_4_op1_tag <= 3'h0; // @[Rob.scala 60:12]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h4 == dispatch_idxs_1) begin // @[Rob.scala 60:12]
        rob_info_4_op1_tag <= 3'h0; // @[Rob.scala 60:12]
      end else begin
        rob_info_4_op1_tag <= _GEN_2980;
      end
    end else begin
      rob_info_4_op1_tag <= _GEN_2980;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_4_op1_data <= 32'h0; // @[Rob.scala 61:13]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_4_op1_data <= 32'h0; // @[Rob.scala 61:13]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h4 == dispatch_idxs_1) begin // @[Rob.scala 61:13]
        rob_info_4_op1_data <= 32'h0; // @[Rob.scala 61:13]
      end else begin
        rob_info_4_op1_data <= _GEN_2988;
      end
    end else begin
      rob_info_4_op1_data <= _GEN_2988;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_4_op2_ready <= 1'h0; // @[Rob.scala 62:14]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_4_op2_ready <= 1'h0; // @[Rob.scala 62:14]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h4 == dispatch_idxs_1) begin // @[Rob.scala 62:14]
        rob_info_4_op2_ready <= 1'h0; // @[Rob.scala 62:14]
      end else begin
        rob_info_4_op2_ready <= _GEN_2996;
      end
    end else begin
      rob_info_4_op2_ready <= _GEN_2996;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_4_op2_tag <= 3'h0; // @[Rob.scala 63:12]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_4_op2_tag <= 3'h0; // @[Rob.scala 63:12]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h4 == dispatch_idxs_1) begin // @[Rob.scala 63:12]
        rob_info_4_op2_tag <= 3'h0; // @[Rob.scala 63:12]
      end else begin
        rob_info_4_op2_tag <= _GEN_3004;
      end
    end else begin
      rob_info_4_op2_tag <= _GEN_3004;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_4_op2_data <= 32'h0; // @[Rob.scala 64:13]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_4_op2_data <= 32'h0; // @[Rob.scala 64:13]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h4 == dispatch_idxs_1) begin // @[Rob.scala 64:13]
        rob_info_4_op2_data <= 32'h0; // @[Rob.scala 64:13]
      end else begin
        rob_info_4_op2_data <= _GEN_3012;
      end
    end else begin
      rob_info_4_op2_data <= _GEN_3012;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_4_imm_data <= 32'h0; // @[Rob.scala 65:13]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_4_imm_data <= 32'h0; // @[Rob.scala 65:13]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h4 == dispatch_idxs_1) begin // @[Rob.scala 65:13]
        rob_info_4_imm_data <= 32'h0; // @[Rob.scala 65:13]
      end else begin
        rob_info_4_imm_data <= _GEN_3020;
      end
    end else begin
      rob_info_4_imm_data <= _GEN_3020;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_4_is_init <= 1'h0; // @[Rob.scala 66:13]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_4_is_init <= 1'h0; // @[Rob.scala 66:13]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h4 == dispatch_idxs_1) begin // @[Rob.scala 66:13]
        rob_info_4_is_init <= 1'h0; // @[Rob.scala 66:13]
      end else begin
        rob_info_4_is_init <= _GEN_3028;
      end
    end else begin
      rob_info_4_is_init <= _GEN_3028;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_4_flush_on_commit <= 1'h0; // @[Rob.scala 67:20]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_4_flush_on_commit <= 1'h0; // @[Rob.scala 67:20]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h4 == dispatch_idxs_1) begin // @[Rob.scala 67:20]
        rob_info_4_flush_on_commit <= 1'h0; // @[Rob.scala 67:20]
      end else begin
        rob_info_4_flush_on_commit <= _GEN_3036;
      end
    end else begin
      rob_info_4_flush_on_commit <= _GEN_3036;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_5_is_valid <= 1'h0; // @[Rob.scala 42:13]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_5_is_valid <= 1'h0; // @[Rob.scala 42:13]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h5 == dispatch_idxs_1) begin // @[Rob.scala 42:13]
        rob_info_5_is_valid <= 1'h0; // @[Rob.scala 42:13]
      end else begin
        rob_info_5_is_valid <= _GEN_2837;
      end
    end else begin
      rob_info_5_is_valid <= _GEN_2837;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_5_busy <= 1'h0; // @[Rob.scala 43:9]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_5_busy <= 1'h0; // @[Rob.scala 43:9]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h5 == dispatch_idxs_1) begin // @[Rob.scala 43:9]
        rob_info_5_busy <= 1'h0; // @[Rob.scala 43:9]
      end else begin
        rob_info_5_busy <= _GEN_2845;
      end
    end else begin
      rob_info_5_busy <= _GEN_2845;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_5_uop <= 6'h0; // @[Rob.scala 44:8]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_5_uop <= 6'h0; // @[Rob.scala 44:8]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h5 == dispatch_idxs_1) begin // @[Rob.scala 44:8]
        rob_info_5_uop <= 6'h0; // @[Rob.scala 44:8]
      end else begin
        rob_info_5_uop <= _GEN_2853;
      end
    end else begin
      rob_info_5_uop <= _GEN_2853;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_5_unit_sel <= 3'h0; // @[Rob.scala 45:13]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_5_unit_sel <= 3'h0; // @[Rob.scala 45:13]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h5 == dispatch_idxs_1) begin // @[Rob.scala 45:13]
        rob_info_5_unit_sel <= 3'h0; // @[Rob.scala 45:13]
      end else begin
        rob_info_5_unit_sel <= _GEN_2861;
      end
    end else begin
      rob_info_5_unit_sel <= _GEN_2861;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_5_need_imm <= 1'h0; // @[Rob.scala 46:13]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_5_need_imm <= 1'h0; // @[Rob.scala 46:13]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h5 == dispatch_idxs_1) begin // @[Rob.scala 46:13]
        rob_info_5_need_imm <= 1'h0; // @[Rob.scala 46:13]
      end else begin
        rob_info_5_need_imm <= _GEN_2869;
      end
    end else begin
      rob_info_5_need_imm <= _GEN_2869;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_5_inst_addr <= 32'h0; // @[Rob.scala 47:14]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_5_inst_addr <= 32'h0; // @[Rob.scala 47:14]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h5 == dispatch_idxs_1) begin // @[Rob.scala 47:14]
        rob_info_5_inst_addr <= 32'h0; // @[Rob.scala 47:14]
      end else begin
        rob_info_5_inst_addr <= _GEN_2877;
      end
    end else begin
      rob_info_5_inst_addr <= _GEN_2877;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_5_commit_addr <= 5'h0; // @[Rob.scala 48:16]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_5_commit_addr <= 5'h0; // @[Rob.scala 48:16]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h5 == dispatch_idxs_1) begin // @[Rob.scala 48:16]
        rob_info_5_commit_addr <= 5'h0; // @[Rob.scala 48:16]
      end else begin
        rob_info_5_commit_addr <= _GEN_2885;
      end
    end else begin
      rob_info_5_commit_addr <= _GEN_2885;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_5_commit_data <= 32'h0; // @[Rob.scala 49:16]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_5_commit_data <= 32'h0; // @[Rob.scala 49:16]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h5 == dispatch_idxs_1) begin // @[Rob.scala 49:16]
        rob_info_5_commit_data <= 32'h0; // @[Rob.scala 49:16]
      end else begin
        rob_info_5_commit_data <= _GEN_2893;
      end
    end else begin
      rob_info_5_commit_data <= _GEN_2893;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_5_commit_ready <= 1'h0; // @[Rob.scala 51:17]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_5_commit_ready <= 1'h0; // @[Rob.scala 51:17]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h5 == dispatch_idxs_1) begin // @[Rob.scala 51:17]
        rob_info_5_commit_ready <= 1'h0; // @[Rob.scala 51:17]
      end else begin
        rob_info_5_commit_ready <= _GEN_2909;
      end
    end else begin
      rob_info_5_commit_ready <= _GEN_2909;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_5_is_branch <= 1'h0; // @[Rob.scala 53:14]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_5_is_branch <= 1'h0; // @[Rob.scala 53:14]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h5 == dispatch_idxs_1) begin // @[Rob.scala 53:14]
        rob_info_5_is_branch <= 1'h0; // @[Rob.scala 53:14]
      end else begin
        rob_info_5_is_branch <= _GEN_2925;
      end
    end else begin
      rob_info_5_is_branch <= _GEN_2925;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_5_predict_taken <= 1'h0; // @[Rob.scala 55:18]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_5_predict_taken <= 1'h0; // @[Rob.scala 55:18]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h5 == dispatch_idxs_1) begin // @[Rob.scala 55:18]
        rob_info_5_predict_taken <= 1'h0; // @[Rob.scala 55:18]
      end else begin
        rob_info_5_predict_taken <= _GEN_2941;
      end
    end else begin
      rob_info_5_predict_taken <= _GEN_2941;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_5_is_taken <= 1'h0; // @[Rob.scala 56:13]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_5_is_taken <= 1'h0; // @[Rob.scala 56:13]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h5 == dispatch_idxs_1) begin // @[Rob.scala 56:13]
        rob_info_5_is_taken <= 1'h0; // @[Rob.scala 56:13]
      end else begin
        rob_info_5_is_taken <= _GEN_2949;
      end
    end else begin
      rob_info_5_is_taken <= _GEN_2949;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_5_predict_miss <= 1'h0; // @[Rob.scala 57:17]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_5_predict_miss <= 1'h0; // @[Rob.scala 57:17]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h5 == dispatch_idxs_1) begin // @[Rob.scala 57:17]
        rob_info_5_predict_miss <= 1'h0; // @[Rob.scala 57:17]
      end else begin
        rob_info_5_predict_miss <= _GEN_2957;
      end
    end else begin
      rob_info_5_predict_miss <= _GEN_2957;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_5_gh_info <= 4'h0; // @[Rob.scala 58:12]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_5_gh_info <= 4'h0; // @[Rob.scala 58:12]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h5 == dispatch_idxs_1) begin // @[Rob.scala 58:12]
        rob_info_5_gh_info <= 4'h0; // @[Rob.scala 58:12]
      end else begin
        rob_info_5_gh_info <= _GEN_2965;
      end
    end else begin
      rob_info_5_gh_info <= _GEN_2965;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_5_op1_ready <= 1'h0; // @[Rob.scala 59:14]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_5_op1_ready <= 1'h0; // @[Rob.scala 59:14]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h5 == dispatch_idxs_1) begin // @[Rob.scala 59:14]
        rob_info_5_op1_ready <= 1'h0; // @[Rob.scala 59:14]
      end else begin
        rob_info_5_op1_ready <= _GEN_2973;
      end
    end else begin
      rob_info_5_op1_ready <= _GEN_2973;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_5_op1_tag <= 3'h0; // @[Rob.scala 60:12]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_5_op1_tag <= 3'h0; // @[Rob.scala 60:12]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h5 == dispatch_idxs_1) begin // @[Rob.scala 60:12]
        rob_info_5_op1_tag <= 3'h0; // @[Rob.scala 60:12]
      end else begin
        rob_info_5_op1_tag <= _GEN_2981;
      end
    end else begin
      rob_info_5_op1_tag <= _GEN_2981;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_5_op1_data <= 32'h0; // @[Rob.scala 61:13]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_5_op1_data <= 32'h0; // @[Rob.scala 61:13]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h5 == dispatch_idxs_1) begin // @[Rob.scala 61:13]
        rob_info_5_op1_data <= 32'h0; // @[Rob.scala 61:13]
      end else begin
        rob_info_5_op1_data <= _GEN_2989;
      end
    end else begin
      rob_info_5_op1_data <= _GEN_2989;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_5_op2_ready <= 1'h0; // @[Rob.scala 62:14]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_5_op2_ready <= 1'h0; // @[Rob.scala 62:14]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h5 == dispatch_idxs_1) begin // @[Rob.scala 62:14]
        rob_info_5_op2_ready <= 1'h0; // @[Rob.scala 62:14]
      end else begin
        rob_info_5_op2_ready <= _GEN_2997;
      end
    end else begin
      rob_info_5_op2_ready <= _GEN_2997;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_5_op2_tag <= 3'h0; // @[Rob.scala 63:12]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_5_op2_tag <= 3'h0; // @[Rob.scala 63:12]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h5 == dispatch_idxs_1) begin // @[Rob.scala 63:12]
        rob_info_5_op2_tag <= 3'h0; // @[Rob.scala 63:12]
      end else begin
        rob_info_5_op2_tag <= _GEN_3005;
      end
    end else begin
      rob_info_5_op2_tag <= _GEN_3005;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_5_op2_data <= 32'h0; // @[Rob.scala 64:13]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_5_op2_data <= 32'h0; // @[Rob.scala 64:13]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h5 == dispatch_idxs_1) begin // @[Rob.scala 64:13]
        rob_info_5_op2_data <= 32'h0; // @[Rob.scala 64:13]
      end else begin
        rob_info_5_op2_data <= _GEN_3013;
      end
    end else begin
      rob_info_5_op2_data <= _GEN_3013;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_5_imm_data <= 32'h0; // @[Rob.scala 65:13]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_5_imm_data <= 32'h0; // @[Rob.scala 65:13]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h5 == dispatch_idxs_1) begin // @[Rob.scala 65:13]
        rob_info_5_imm_data <= 32'h0; // @[Rob.scala 65:13]
      end else begin
        rob_info_5_imm_data <= _GEN_3021;
      end
    end else begin
      rob_info_5_imm_data <= _GEN_3021;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_5_is_init <= 1'h0; // @[Rob.scala 66:13]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_5_is_init <= 1'h0; // @[Rob.scala 66:13]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h5 == dispatch_idxs_1) begin // @[Rob.scala 66:13]
        rob_info_5_is_init <= 1'h0; // @[Rob.scala 66:13]
      end else begin
        rob_info_5_is_init <= _GEN_3029;
      end
    end else begin
      rob_info_5_is_init <= _GEN_3029;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_5_flush_on_commit <= 1'h0; // @[Rob.scala 67:20]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_5_flush_on_commit <= 1'h0; // @[Rob.scala 67:20]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h5 == dispatch_idxs_1) begin // @[Rob.scala 67:20]
        rob_info_5_flush_on_commit <= 1'h0; // @[Rob.scala 67:20]
      end else begin
        rob_info_5_flush_on_commit <= _GEN_3037;
      end
    end else begin
      rob_info_5_flush_on_commit <= _GEN_3037;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_6_is_valid <= 1'h0; // @[Rob.scala 42:13]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_6_is_valid <= 1'h0; // @[Rob.scala 42:13]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h6 == dispatch_idxs_1) begin // @[Rob.scala 42:13]
        rob_info_6_is_valid <= 1'h0; // @[Rob.scala 42:13]
      end else begin
        rob_info_6_is_valid <= _GEN_2838;
      end
    end else begin
      rob_info_6_is_valid <= _GEN_2838;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_6_busy <= 1'h0; // @[Rob.scala 43:9]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_6_busy <= 1'h0; // @[Rob.scala 43:9]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h6 == dispatch_idxs_1) begin // @[Rob.scala 43:9]
        rob_info_6_busy <= 1'h0; // @[Rob.scala 43:9]
      end else begin
        rob_info_6_busy <= _GEN_2846;
      end
    end else begin
      rob_info_6_busy <= _GEN_2846;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_6_uop <= 6'h0; // @[Rob.scala 44:8]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_6_uop <= 6'h0; // @[Rob.scala 44:8]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h6 == dispatch_idxs_1) begin // @[Rob.scala 44:8]
        rob_info_6_uop <= 6'h0; // @[Rob.scala 44:8]
      end else begin
        rob_info_6_uop <= _GEN_2854;
      end
    end else begin
      rob_info_6_uop <= _GEN_2854;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_6_unit_sel <= 3'h0; // @[Rob.scala 45:13]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_6_unit_sel <= 3'h0; // @[Rob.scala 45:13]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h6 == dispatch_idxs_1) begin // @[Rob.scala 45:13]
        rob_info_6_unit_sel <= 3'h0; // @[Rob.scala 45:13]
      end else begin
        rob_info_6_unit_sel <= _GEN_2862;
      end
    end else begin
      rob_info_6_unit_sel <= _GEN_2862;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_6_need_imm <= 1'h0; // @[Rob.scala 46:13]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_6_need_imm <= 1'h0; // @[Rob.scala 46:13]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h6 == dispatch_idxs_1) begin // @[Rob.scala 46:13]
        rob_info_6_need_imm <= 1'h0; // @[Rob.scala 46:13]
      end else begin
        rob_info_6_need_imm <= _GEN_2870;
      end
    end else begin
      rob_info_6_need_imm <= _GEN_2870;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_6_inst_addr <= 32'h0; // @[Rob.scala 47:14]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_6_inst_addr <= 32'h0; // @[Rob.scala 47:14]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h6 == dispatch_idxs_1) begin // @[Rob.scala 47:14]
        rob_info_6_inst_addr <= 32'h0; // @[Rob.scala 47:14]
      end else begin
        rob_info_6_inst_addr <= _GEN_2878;
      end
    end else begin
      rob_info_6_inst_addr <= _GEN_2878;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_6_commit_addr <= 5'h0; // @[Rob.scala 48:16]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_6_commit_addr <= 5'h0; // @[Rob.scala 48:16]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h6 == dispatch_idxs_1) begin // @[Rob.scala 48:16]
        rob_info_6_commit_addr <= 5'h0; // @[Rob.scala 48:16]
      end else begin
        rob_info_6_commit_addr <= _GEN_2886;
      end
    end else begin
      rob_info_6_commit_addr <= _GEN_2886;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_6_commit_data <= 32'h0; // @[Rob.scala 49:16]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_6_commit_data <= 32'h0; // @[Rob.scala 49:16]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h6 == dispatch_idxs_1) begin // @[Rob.scala 49:16]
        rob_info_6_commit_data <= 32'h0; // @[Rob.scala 49:16]
      end else begin
        rob_info_6_commit_data <= _GEN_2894;
      end
    end else begin
      rob_info_6_commit_data <= _GEN_2894;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_6_commit_ready <= 1'h0; // @[Rob.scala 51:17]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_6_commit_ready <= 1'h0; // @[Rob.scala 51:17]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h6 == dispatch_idxs_1) begin // @[Rob.scala 51:17]
        rob_info_6_commit_ready <= 1'h0; // @[Rob.scala 51:17]
      end else begin
        rob_info_6_commit_ready <= _GEN_2910;
      end
    end else begin
      rob_info_6_commit_ready <= _GEN_2910;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_6_is_branch <= 1'h0; // @[Rob.scala 53:14]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_6_is_branch <= 1'h0; // @[Rob.scala 53:14]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h6 == dispatch_idxs_1) begin // @[Rob.scala 53:14]
        rob_info_6_is_branch <= 1'h0; // @[Rob.scala 53:14]
      end else begin
        rob_info_6_is_branch <= _GEN_2926;
      end
    end else begin
      rob_info_6_is_branch <= _GEN_2926;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_6_predict_taken <= 1'h0; // @[Rob.scala 55:18]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_6_predict_taken <= 1'h0; // @[Rob.scala 55:18]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h6 == dispatch_idxs_1) begin // @[Rob.scala 55:18]
        rob_info_6_predict_taken <= 1'h0; // @[Rob.scala 55:18]
      end else begin
        rob_info_6_predict_taken <= _GEN_2942;
      end
    end else begin
      rob_info_6_predict_taken <= _GEN_2942;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_6_is_taken <= 1'h0; // @[Rob.scala 56:13]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_6_is_taken <= 1'h0; // @[Rob.scala 56:13]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h6 == dispatch_idxs_1) begin // @[Rob.scala 56:13]
        rob_info_6_is_taken <= 1'h0; // @[Rob.scala 56:13]
      end else begin
        rob_info_6_is_taken <= _GEN_2950;
      end
    end else begin
      rob_info_6_is_taken <= _GEN_2950;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_6_predict_miss <= 1'h0; // @[Rob.scala 57:17]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_6_predict_miss <= 1'h0; // @[Rob.scala 57:17]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h6 == dispatch_idxs_1) begin // @[Rob.scala 57:17]
        rob_info_6_predict_miss <= 1'h0; // @[Rob.scala 57:17]
      end else begin
        rob_info_6_predict_miss <= _GEN_2958;
      end
    end else begin
      rob_info_6_predict_miss <= _GEN_2958;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_6_gh_info <= 4'h0; // @[Rob.scala 58:12]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_6_gh_info <= 4'h0; // @[Rob.scala 58:12]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h6 == dispatch_idxs_1) begin // @[Rob.scala 58:12]
        rob_info_6_gh_info <= 4'h0; // @[Rob.scala 58:12]
      end else begin
        rob_info_6_gh_info <= _GEN_2966;
      end
    end else begin
      rob_info_6_gh_info <= _GEN_2966;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_6_op1_ready <= 1'h0; // @[Rob.scala 59:14]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_6_op1_ready <= 1'h0; // @[Rob.scala 59:14]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h6 == dispatch_idxs_1) begin // @[Rob.scala 59:14]
        rob_info_6_op1_ready <= 1'h0; // @[Rob.scala 59:14]
      end else begin
        rob_info_6_op1_ready <= _GEN_2974;
      end
    end else begin
      rob_info_6_op1_ready <= _GEN_2974;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_6_op1_tag <= 3'h0; // @[Rob.scala 60:12]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_6_op1_tag <= 3'h0; // @[Rob.scala 60:12]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h6 == dispatch_idxs_1) begin // @[Rob.scala 60:12]
        rob_info_6_op1_tag <= 3'h0; // @[Rob.scala 60:12]
      end else begin
        rob_info_6_op1_tag <= _GEN_2982;
      end
    end else begin
      rob_info_6_op1_tag <= _GEN_2982;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_6_op1_data <= 32'h0; // @[Rob.scala 61:13]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_6_op1_data <= 32'h0; // @[Rob.scala 61:13]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h6 == dispatch_idxs_1) begin // @[Rob.scala 61:13]
        rob_info_6_op1_data <= 32'h0; // @[Rob.scala 61:13]
      end else begin
        rob_info_6_op1_data <= _GEN_2990;
      end
    end else begin
      rob_info_6_op1_data <= _GEN_2990;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_6_op2_ready <= 1'h0; // @[Rob.scala 62:14]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_6_op2_ready <= 1'h0; // @[Rob.scala 62:14]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h6 == dispatch_idxs_1) begin // @[Rob.scala 62:14]
        rob_info_6_op2_ready <= 1'h0; // @[Rob.scala 62:14]
      end else begin
        rob_info_6_op2_ready <= _GEN_2998;
      end
    end else begin
      rob_info_6_op2_ready <= _GEN_2998;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_6_op2_tag <= 3'h0; // @[Rob.scala 63:12]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_6_op2_tag <= 3'h0; // @[Rob.scala 63:12]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h6 == dispatch_idxs_1) begin // @[Rob.scala 63:12]
        rob_info_6_op2_tag <= 3'h0; // @[Rob.scala 63:12]
      end else begin
        rob_info_6_op2_tag <= _GEN_3006;
      end
    end else begin
      rob_info_6_op2_tag <= _GEN_3006;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_6_op2_data <= 32'h0; // @[Rob.scala 64:13]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_6_op2_data <= 32'h0; // @[Rob.scala 64:13]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h6 == dispatch_idxs_1) begin // @[Rob.scala 64:13]
        rob_info_6_op2_data <= 32'h0; // @[Rob.scala 64:13]
      end else begin
        rob_info_6_op2_data <= _GEN_3014;
      end
    end else begin
      rob_info_6_op2_data <= _GEN_3014;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_6_imm_data <= 32'h0; // @[Rob.scala 65:13]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_6_imm_data <= 32'h0; // @[Rob.scala 65:13]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h6 == dispatch_idxs_1) begin // @[Rob.scala 65:13]
        rob_info_6_imm_data <= 32'h0; // @[Rob.scala 65:13]
      end else begin
        rob_info_6_imm_data <= _GEN_3022;
      end
    end else begin
      rob_info_6_imm_data <= _GEN_3022;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_6_is_init <= 1'h0; // @[Rob.scala 66:13]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_6_is_init <= 1'h0; // @[Rob.scala 66:13]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h6 == dispatch_idxs_1) begin // @[Rob.scala 66:13]
        rob_info_6_is_init <= 1'h0; // @[Rob.scala 66:13]
      end else begin
        rob_info_6_is_init <= _GEN_3030;
      end
    end else begin
      rob_info_6_is_init <= _GEN_3030;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_6_flush_on_commit <= 1'h0; // @[Rob.scala 67:20]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_6_flush_on_commit <= 1'h0; // @[Rob.scala 67:20]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h6 == dispatch_idxs_1) begin // @[Rob.scala 67:20]
        rob_info_6_flush_on_commit <= 1'h0; // @[Rob.scala 67:20]
      end else begin
        rob_info_6_flush_on_commit <= _GEN_3038;
      end
    end else begin
      rob_info_6_flush_on_commit <= _GEN_3038;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_7_is_valid <= 1'h0; // @[Rob.scala 42:13]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_7_is_valid <= 1'h0; // @[Rob.scala 42:13]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h7 == dispatch_idxs_1) begin // @[Rob.scala 42:13]
        rob_info_7_is_valid <= 1'h0; // @[Rob.scala 42:13]
      end else begin
        rob_info_7_is_valid <= _GEN_2839;
      end
    end else begin
      rob_info_7_is_valid <= _GEN_2839;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_7_busy <= 1'h0; // @[Rob.scala 43:9]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_7_busy <= 1'h0; // @[Rob.scala 43:9]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h7 == dispatch_idxs_1) begin // @[Rob.scala 43:9]
        rob_info_7_busy <= 1'h0; // @[Rob.scala 43:9]
      end else begin
        rob_info_7_busy <= _GEN_2847;
      end
    end else begin
      rob_info_7_busy <= _GEN_2847;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_7_uop <= 6'h0; // @[Rob.scala 44:8]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_7_uop <= 6'h0; // @[Rob.scala 44:8]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h7 == dispatch_idxs_1) begin // @[Rob.scala 44:8]
        rob_info_7_uop <= 6'h0; // @[Rob.scala 44:8]
      end else begin
        rob_info_7_uop <= _GEN_2855;
      end
    end else begin
      rob_info_7_uop <= _GEN_2855;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_7_unit_sel <= 3'h0; // @[Rob.scala 45:13]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_7_unit_sel <= 3'h0; // @[Rob.scala 45:13]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h7 == dispatch_idxs_1) begin // @[Rob.scala 45:13]
        rob_info_7_unit_sel <= 3'h0; // @[Rob.scala 45:13]
      end else begin
        rob_info_7_unit_sel <= _GEN_2863;
      end
    end else begin
      rob_info_7_unit_sel <= _GEN_2863;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_7_need_imm <= 1'h0; // @[Rob.scala 46:13]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_7_need_imm <= 1'h0; // @[Rob.scala 46:13]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h7 == dispatch_idxs_1) begin // @[Rob.scala 46:13]
        rob_info_7_need_imm <= 1'h0; // @[Rob.scala 46:13]
      end else begin
        rob_info_7_need_imm <= _GEN_2871;
      end
    end else begin
      rob_info_7_need_imm <= _GEN_2871;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_7_inst_addr <= 32'h0; // @[Rob.scala 47:14]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_7_inst_addr <= 32'h0; // @[Rob.scala 47:14]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h7 == dispatch_idxs_1) begin // @[Rob.scala 47:14]
        rob_info_7_inst_addr <= 32'h0; // @[Rob.scala 47:14]
      end else begin
        rob_info_7_inst_addr <= _GEN_2879;
      end
    end else begin
      rob_info_7_inst_addr <= _GEN_2879;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_7_commit_addr <= 5'h0; // @[Rob.scala 48:16]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_7_commit_addr <= 5'h0; // @[Rob.scala 48:16]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h7 == dispatch_idxs_1) begin // @[Rob.scala 48:16]
        rob_info_7_commit_addr <= 5'h0; // @[Rob.scala 48:16]
      end else begin
        rob_info_7_commit_addr <= _GEN_2887;
      end
    end else begin
      rob_info_7_commit_addr <= _GEN_2887;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_7_commit_data <= 32'h0; // @[Rob.scala 49:16]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_7_commit_data <= 32'h0; // @[Rob.scala 49:16]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h7 == dispatch_idxs_1) begin // @[Rob.scala 49:16]
        rob_info_7_commit_data <= 32'h0; // @[Rob.scala 49:16]
      end else begin
        rob_info_7_commit_data <= _GEN_2895;
      end
    end else begin
      rob_info_7_commit_data <= _GEN_2895;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_7_commit_ready <= 1'h0; // @[Rob.scala 51:17]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_7_commit_ready <= 1'h0; // @[Rob.scala 51:17]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h7 == dispatch_idxs_1) begin // @[Rob.scala 51:17]
        rob_info_7_commit_ready <= 1'h0; // @[Rob.scala 51:17]
      end else begin
        rob_info_7_commit_ready <= _GEN_2911;
      end
    end else begin
      rob_info_7_commit_ready <= _GEN_2911;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_7_is_branch <= 1'h0; // @[Rob.scala 53:14]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_7_is_branch <= 1'h0; // @[Rob.scala 53:14]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h7 == dispatch_idxs_1) begin // @[Rob.scala 53:14]
        rob_info_7_is_branch <= 1'h0; // @[Rob.scala 53:14]
      end else begin
        rob_info_7_is_branch <= _GEN_2927;
      end
    end else begin
      rob_info_7_is_branch <= _GEN_2927;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_7_predict_taken <= 1'h0; // @[Rob.scala 55:18]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_7_predict_taken <= 1'h0; // @[Rob.scala 55:18]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h7 == dispatch_idxs_1) begin // @[Rob.scala 55:18]
        rob_info_7_predict_taken <= 1'h0; // @[Rob.scala 55:18]
      end else begin
        rob_info_7_predict_taken <= _GEN_2943;
      end
    end else begin
      rob_info_7_predict_taken <= _GEN_2943;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_7_is_taken <= 1'h0; // @[Rob.scala 56:13]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_7_is_taken <= 1'h0; // @[Rob.scala 56:13]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h7 == dispatch_idxs_1) begin // @[Rob.scala 56:13]
        rob_info_7_is_taken <= 1'h0; // @[Rob.scala 56:13]
      end else begin
        rob_info_7_is_taken <= _GEN_2951;
      end
    end else begin
      rob_info_7_is_taken <= _GEN_2951;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_7_predict_miss <= 1'h0; // @[Rob.scala 57:17]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_7_predict_miss <= 1'h0; // @[Rob.scala 57:17]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h7 == dispatch_idxs_1) begin // @[Rob.scala 57:17]
        rob_info_7_predict_miss <= 1'h0; // @[Rob.scala 57:17]
      end else begin
        rob_info_7_predict_miss <= _GEN_2959;
      end
    end else begin
      rob_info_7_predict_miss <= _GEN_2959;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_7_gh_info <= 4'h0; // @[Rob.scala 58:12]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_7_gh_info <= 4'h0; // @[Rob.scala 58:12]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h7 == dispatch_idxs_1) begin // @[Rob.scala 58:12]
        rob_info_7_gh_info <= 4'h0; // @[Rob.scala 58:12]
      end else begin
        rob_info_7_gh_info <= _GEN_2967;
      end
    end else begin
      rob_info_7_gh_info <= _GEN_2967;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_7_op1_ready <= 1'h0; // @[Rob.scala 59:14]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_7_op1_ready <= 1'h0; // @[Rob.scala 59:14]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h7 == dispatch_idxs_1) begin // @[Rob.scala 59:14]
        rob_info_7_op1_ready <= 1'h0; // @[Rob.scala 59:14]
      end else begin
        rob_info_7_op1_ready <= _GEN_2975;
      end
    end else begin
      rob_info_7_op1_ready <= _GEN_2975;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_7_op1_tag <= 3'h0; // @[Rob.scala 60:12]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_7_op1_tag <= 3'h0; // @[Rob.scala 60:12]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h7 == dispatch_idxs_1) begin // @[Rob.scala 60:12]
        rob_info_7_op1_tag <= 3'h0; // @[Rob.scala 60:12]
      end else begin
        rob_info_7_op1_tag <= _GEN_2983;
      end
    end else begin
      rob_info_7_op1_tag <= _GEN_2983;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_7_op1_data <= 32'h0; // @[Rob.scala 61:13]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_7_op1_data <= 32'h0; // @[Rob.scala 61:13]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h7 == dispatch_idxs_1) begin // @[Rob.scala 61:13]
        rob_info_7_op1_data <= 32'h0; // @[Rob.scala 61:13]
      end else begin
        rob_info_7_op1_data <= _GEN_2991;
      end
    end else begin
      rob_info_7_op1_data <= _GEN_2991;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_7_op2_ready <= 1'h0; // @[Rob.scala 62:14]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_7_op2_ready <= 1'h0; // @[Rob.scala 62:14]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h7 == dispatch_idxs_1) begin // @[Rob.scala 62:14]
        rob_info_7_op2_ready <= 1'h0; // @[Rob.scala 62:14]
      end else begin
        rob_info_7_op2_ready <= _GEN_2999;
      end
    end else begin
      rob_info_7_op2_ready <= _GEN_2999;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_7_op2_tag <= 3'h0; // @[Rob.scala 63:12]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_7_op2_tag <= 3'h0; // @[Rob.scala 63:12]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h7 == dispatch_idxs_1) begin // @[Rob.scala 63:12]
        rob_info_7_op2_tag <= 3'h0; // @[Rob.scala 63:12]
      end else begin
        rob_info_7_op2_tag <= _GEN_3007;
      end
    end else begin
      rob_info_7_op2_tag <= _GEN_3007;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_7_op2_data <= 32'h0; // @[Rob.scala 64:13]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_7_op2_data <= 32'h0; // @[Rob.scala 64:13]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h7 == dispatch_idxs_1) begin // @[Rob.scala 64:13]
        rob_info_7_op2_data <= 32'h0; // @[Rob.scala 64:13]
      end else begin
        rob_info_7_op2_data <= _GEN_3015;
      end
    end else begin
      rob_info_7_op2_data <= _GEN_3015;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_7_imm_data <= 32'h0; // @[Rob.scala 65:13]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_7_imm_data <= 32'h0; // @[Rob.scala 65:13]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h7 == dispatch_idxs_1) begin // @[Rob.scala 65:13]
        rob_info_7_imm_data <= 32'h0; // @[Rob.scala 65:13]
      end else begin
        rob_info_7_imm_data <= _GEN_3023;
      end
    end else begin
      rob_info_7_imm_data <= _GEN_3023;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_7_is_init <= 1'h0; // @[Rob.scala 66:13]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_7_is_init <= 1'h0; // @[Rob.scala 66:13]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h7 == dispatch_idxs_1) begin // @[Rob.scala 66:13]
        rob_info_7_is_init <= 1'h0; // @[Rob.scala 66:13]
      end else begin
        rob_info_7_is_init <= _GEN_3031;
      end
    end else begin
      rob_info_7_is_init <= _GEN_3031;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_info_7_flush_on_commit <= 1'h0; // @[Rob.scala 67:20]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_info_7_flush_on_commit <= 1'h0; // @[Rob.scala 67:20]
    end else if (deq_ready_mask_1) begin // @[Rob.scala 349:28]
      if (3'h7 == dispatch_idxs_1) begin // @[Rob.scala 67:20]
        rob_info_7_flush_on_commit <= 1'h0; // @[Rob.scala 67:20]
      end else begin
        rob_info_7_flush_on_commit <= _GEN_3039;
      end
    end else begin
      rob_info_7_flush_on_commit <= _GEN_3039;
    end
    if (reset) begin // @[Rob.scala 176:31]
      head <= 8'h1; // @[Rob.scala 176:31]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      head <= _dispatch_idxs_T_3; // @[Rob.scala 459:10]
    end else if (2'h2 == _head_next_T_1) begin // @[Rob.scala 333:20]
      head <= _dispatch_idxs_T_7; // @[Rob.scala 333:20]
    end else if (2'h1 == _head_next_T_1) begin // @[Rob.scala 333:20]
      head <= _dispatch_idxs_T_3; // @[Rob.scala 333:20]
    end
    if (reset) begin // @[Rob.scala 178:31]
      tail <= 8'h1; // @[Rob.scala 178:31]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      tail <= _dispatch_idxs_T_3; // @[Rob.scala 458:10]
    end else if (inst_valid_mask_1 & ~might_hit_1) begin // @[Rob.scala 195:20]
      tail <= _T_13;
    end else if (inst_valid_mask_0 & ~might_hit_head_mask_0) begin // @[Rob.scala 195:20]
      tail <= _T_6;
    end
    if (reset) begin // @[Rob.scala 179:31]
      maybe_full <= 1'h0; // @[Rob.scala 179:31]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      maybe_full <= 1'h0; // @[Rob.scala 460:16]
    end else begin
      maybe_full <= _GEN_3579;
    end
    if (reset) begin // @[Rob.scala 187:30]
      waiting_delay <= 1'h0; // @[Rob.scala 187:30]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      waiting_delay <= 1'h0; // @[Rob.scala 461:18]
    end else if (waiting_delay) begin // @[Rob.scala 429:22]
      if (deq_ready_mask_0) begin // @[Rob.scala 432:28]
        waiting_delay <= 1'h0; // @[Rob.scala 433:20]
      end else begin
        waiting_delay <= _GEN_3580;
      end
    end else begin
      waiting_delay <= _GEN_3580;
    end
    if (reset) begin // @[Rob.scala 188:27]
      need_flush <= 1'h0; // @[Rob.scala 188:27]
    end else begin
      need_flush <= _GEN_3591;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_commit_1_des_rob <= 3'h0; // @[Rename.scala 15:13]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_commit_1_des_rob <= 3'h0; // @[Rename.scala 15:13]
    end else begin
      rob_commit_1_des_rob <= dispatch_idxs_1; // @[Rob.scala 347:27]
    end
    if (reset) begin // @[Rob.scala 342:33]
      rob_commit_valid_1 <= 1'h0; // @[Rob.scala 342:33]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_commit_valid_1 <= 1'h0; // @[Rob.scala 456:8]
    end else if (waiting_delay) begin // @[Rob.scala 429:22]
      rob_commit_valid_1 <= 1'h0; // @[Rob.scala 430:58]
    end else begin
      rob_commit_valid_1 <= deq_ready_mask_1; // @[Rob.scala 345:25]
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_commit_0_des_rob <= 3'h0; // @[Rename.scala 15:13]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_commit_0_des_rob <= 3'h0; // @[Rename.scala 15:13]
    end else begin
      rob_commit_0_des_rob <= dispatch_idxs_0; // @[Rob.scala 347:27]
    end
    if (reset) begin // @[Rob.scala 342:33]
      rob_commit_valid_0 <= 1'h0; // @[Rob.scala 342:33]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_commit_valid_0 <= 1'h0; // @[Rob.scala 456:8]
    end else begin
      rob_commit_valid_0 <= deq_ready_mask_0; // @[Rob.scala 345:25]
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_commit_1_commit_data <= 32'h0; // @[Rename.scala 17:17]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_commit_1_commit_data <= 32'h0; // @[Rename.scala 17:17]
    end else if (3'h7 == dispatch_idxs_1) begin // @[Rob.scala 346:31]
      rob_commit_1_commit_data <= rob_info_7_commit_data; // @[Rob.scala 346:31]
    end else if (3'h6 == dispatch_idxs_1) begin // @[Rob.scala 346:31]
      rob_commit_1_commit_data <= rob_info_6_commit_data; // @[Rob.scala 346:31]
    end else begin
      rob_commit_1_commit_data <= _GEN_3045;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_commit_0_commit_data <= 32'h0; // @[Rename.scala 17:17]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_commit_0_commit_data <= 32'h0; // @[Rename.scala 17:17]
    end else if (3'h7 == dispatch_idxs_0) begin // @[Rob.scala 346:31]
      rob_commit_0_commit_data <= rob_info_7_commit_data; // @[Rob.scala 346:31]
    end else if (3'h6 == dispatch_idxs_0) begin // @[Rob.scala 346:31]
      rob_commit_0_commit_data <= rob_info_6_commit_data; // @[Rob.scala 346:31]
    end else begin
      rob_commit_0_commit_data <= _GEN_2613;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_commit_0_commit_addr <= 5'h0; // @[Rename.scala 16:17]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_commit_0_commit_addr <= 5'h0; // @[Rename.scala 16:17]
    end else if (3'h7 == dispatch_idxs_0) begin // @[Rob.scala 348:31]
      rob_commit_0_commit_addr <= rob_info_7_commit_addr; // @[Rob.scala 348:31]
    end else if (3'h6 == dispatch_idxs_0) begin // @[Rob.scala 348:31]
      rob_commit_0_commit_addr <= rob_info_6_commit_addr; // @[Rob.scala 348:31]
    end else begin
      rob_commit_0_commit_addr <= _GEN_2621;
    end
    if (reset) begin // @[Rob.scala 464:24]
      rob_commit_1_commit_addr <= 5'h0; // @[Rename.scala 16:17]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      rob_commit_1_commit_addr <= 5'h0; // @[Rename.scala 16:17]
    end else if (3'h7 == dispatch_idxs_1) begin // @[Rob.scala 348:31]
      rob_commit_1_commit_addr <= rob_info_7_commit_addr; // @[Rob.scala 348:31]
    end else if (3'h6 == dispatch_idxs_1) begin // @[Rob.scala 348:31]
      rob_commit_1_commit_addr <= rob_info_6_commit_addr; // @[Rob.scala 348:31]
    end else begin
      rob_commit_1_commit_addr <= _GEN_3053;
    end
    if (reset) begin // @[Rob.scala 464:24]
      branch_info_target_addr <= 32'h0; // @[Bpu.scala 42:18]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      branch_info_target_addr <= 32'h0; // @[Bpu.scala 42:18]
    end else if (!(waiting_delay)) begin // @[Rob.scala 429:22]
      if (3'h7 == _GEN_3529) begin // @[Rob.scala 388:27]
        branch_info_target_addr <= rob_info_7_imm_data; // @[Rob.scala 388:27]
      end else begin
        branch_info_target_addr <= _GEN_3536;
      end
    end
    if (reset) begin // @[Rob.scala 464:24]
      branch_info_inst_addr <= 32'h0; // @[Bpu.scala 43:18]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      branch_info_inst_addr <= 32'h0; // @[Bpu.scala 43:18]
    end else if (!(waiting_delay)) begin // @[Rob.scala 429:22]
      if (3'h7 == _GEN_3529) begin // @[Rob.scala 389:25]
        branch_info_inst_addr <= rob_info_7_inst_addr; // @[Rob.scala 389:25]
      end else begin
        branch_info_inst_addr <= _GEN_3544;
      end
    end
    if (reset) begin // @[Rob.scala 464:24]
      branch_info_gh_update <= 4'h0; // @[Bpu.scala 44:18]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      branch_info_gh_update <= 4'h0; // @[Bpu.scala 44:18]
    end else if (!(waiting_delay)) begin // @[Rob.scala 429:22]
      if (3'h7 == _GEN_3529) begin // @[Rob.scala 390:25]
        branch_info_gh_update <= rob_info_7_gh_info; // @[Rob.scala 390:25]
      end else begin
        branch_info_gh_update <= _GEN_3552;
      end
    end
    if (reset) begin // @[Rob.scala 464:24]
      branch_info_is_branch <= 1'h0; // @[Bpu.scala 45:18]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      branch_info_is_branch <= 1'h0; // @[Bpu.scala 45:18]
    end else if (!(waiting_delay)) begin // @[Rob.scala 429:22]
      if (3'h7 == _GEN_3529) begin // @[Rob.scala 391:25]
        branch_info_is_branch <= rob_info_7_is_branch; // @[Rob.scala 391:25]
      end else begin
        branch_info_is_branch <= _GEN_3560;
      end
    end
    if (reset) begin // @[Rob.scala 464:24]
      branch_info_is_taken <= 1'h0; // @[Bpu.scala 46:18]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      branch_info_is_taken <= 1'h0; // @[Bpu.scala 46:18]
    end else if (!(waiting_delay)) begin // @[Rob.scala 429:22]
      if (3'h7 == _GEN_3529) begin // @[Rob.scala 392:24]
        branch_info_is_taken <= rob_info_7_is_taken; // @[Rob.scala 392:24]
      end else begin
        branch_info_is_taken <= _GEN_3568;
      end
    end
    if (reset) begin // @[Rob.scala 464:24]
      branch_info_predict_miss <= 1'h0; // @[Bpu.scala 47:18]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      branch_info_predict_miss <= 1'h0; // @[Bpu.scala 47:18]
    end else if (!(waiting_delay)) begin // @[Rob.scala 429:22]
      if (3'h7 == _GEN_3529) begin // @[Rob.scala 393:28]
        branch_info_predict_miss <= rob_info_7_predict_miss; // @[Rob.scala 393:28]
      end else begin
        branch_info_predict_miss <= _GEN_3576;
      end
    end
    if (reset) begin // @[Rob.scala 386:34]
      branch_info_valid <= 1'h0; // @[Rob.scala 386:34]
    end else if (need_flush) begin // @[Rob.scala 445:19]
      branch_info_valid <= 1'h0; // @[Rob.scala 450:22]
    end else begin
      branch_info_valid <= _GEN_3591;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  rob_info_0_is_valid = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  rob_info_0_busy = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  rob_info_0_uop = _RAND_2[5:0];
  _RAND_3 = {1{`RANDOM}};
  rob_info_0_unit_sel = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  rob_info_0_need_imm = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  rob_info_0_inst_addr = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  rob_info_0_commit_addr = _RAND_6[4:0];
  _RAND_7 = {1{`RANDOM}};
  rob_info_0_commit_data = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  rob_info_0_commit_ready = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  rob_info_0_is_branch = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  rob_info_0_predict_taken = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  rob_info_0_is_taken = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  rob_info_0_predict_miss = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  rob_info_0_gh_info = _RAND_13[3:0];
  _RAND_14 = {1{`RANDOM}};
  rob_info_0_op1_ready = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  rob_info_0_op1_tag = _RAND_15[2:0];
  _RAND_16 = {1{`RANDOM}};
  rob_info_0_op1_data = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  rob_info_0_op2_ready = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  rob_info_0_op2_tag = _RAND_18[2:0];
  _RAND_19 = {1{`RANDOM}};
  rob_info_0_op2_data = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  rob_info_0_imm_data = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  rob_info_0_is_init = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  rob_info_0_flush_on_commit = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  rob_info_1_is_valid = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  rob_info_1_busy = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  rob_info_1_uop = _RAND_25[5:0];
  _RAND_26 = {1{`RANDOM}};
  rob_info_1_unit_sel = _RAND_26[2:0];
  _RAND_27 = {1{`RANDOM}};
  rob_info_1_need_imm = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  rob_info_1_inst_addr = _RAND_28[31:0];
  _RAND_29 = {1{`RANDOM}};
  rob_info_1_commit_addr = _RAND_29[4:0];
  _RAND_30 = {1{`RANDOM}};
  rob_info_1_commit_data = _RAND_30[31:0];
  _RAND_31 = {1{`RANDOM}};
  rob_info_1_commit_ready = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  rob_info_1_is_branch = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  rob_info_1_predict_taken = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  rob_info_1_is_taken = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  rob_info_1_predict_miss = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  rob_info_1_gh_info = _RAND_36[3:0];
  _RAND_37 = {1{`RANDOM}};
  rob_info_1_op1_ready = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  rob_info_1_op1_tag = _RAND_38[2:0];
  _RAND_39 = {1{`RANDOM}};
  rob_info_1_op1_data = _RAND_39[31:0];
  _RAND_40 = {1{`RANDOM}};
  rob_info_1_op2_ready = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  rob_info_1_op2_tag = _RAND_41[2:0];
  _RAND_42 = {1{`RANDOM}};
  rob_info_1_op2_data = _RAND_42[31:0];
  _RAND_43 = {1{`RANDOM}};
  rob_info_1_imm_data = _RAND_43[31:0];
  _RAND_44 = {1{`RANDOM}};
  rob_info_1_is_init = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  rob_info_1_flush_on_commit = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  rob_info_2_is_valid = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  rob_info_2_busy = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  rob_info_2_uop = _RAND_48[5:0];
  _RAND_49 = {1{`RANDOM}};
  rob_info_2_unit_sel = _RAND_49[2:0];
  _RAND_50 = {1{`RANDOM}};
  rob_info_2_need_imm = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  rob_info_2_inst_addr = _RAND_51[31:0];
  _RAND_52 = {1{`RANDOM}};
  rob_info_2_commit_addr = _RAND_52[4:0];
  _RAND_53 = {1{`RANDOM}};
  rob_info_2_commit_data = _RAND_53[31:0];
  _RAND_54 = {1{`RANDOM}};
  rob_info_2_commit_ready = _RAND_54[0:0];
  _RAND_55 = {1{`RANDOM}};
  rob_info_2_is_branch = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  rob_info_2_predict_taken = _RAND_56[0:0];
  _RAND_57 = {1{`RANDOM}};
  rob_info_2_is_taken = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  rob_info_2_predict_miss = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  rob_info_2_gh_info = _RAND_59[3:0];
  _RAND_60 = {1{`RANDOM}};
  rob_info_2_op1_ready = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  rob_info_2_op1_tag = _RAND_61[2:0];
  _RAND_62 = {1{`RANDOM}};
  rob_info_2_op1_data = _RAND_62[31:0];
  _RAND_63 = {1{`RANDOM}};
  rob_info_2_op2_ready = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  rob_info_2_op2_tag = _RAND_64[2:0];
  _RAND_65 = {1{`RANDOM}};
  rob_info_2_op2_data = _RAND_65[31:0];
  _RAND_66 = {1{`RANDOM}};
  rob_info_2_imm_data = _RAND_66[31:0];
  _RAND_67 = {1{`RANDOM}};
  rob_info_2_is_init = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  rob_info_2_flush_on_commit = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  rob_info_3_is_valid = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  rob_info_3_busy = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  rob_info_3_uop = _RAND_71[5:0];
  _RAND_72 = {1{`RANDOM}};
  rob_info_3_unit_sel = _RAND_72[2:0];
  _RAND_73 = {1{`RANDOM}};
  rob_info_3_need_imm = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  rob_info_3_inst_addr = _RAND_74[31:0];
  _RAND_75 = {1{`RANDOM}};
  rob_info_3_commit_addr = _RAND_75[4:0];
  _RAND_76 = {1{`RANDOM}};
  rob_info_3_commit_data = _RAND_76[31:0];
  _RAND_77 = {1{`RANDOM}};
  rob_info_3_commit_ready = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  rob_info_3_is_branch = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  rob_info_3_predict_taken = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  rob_info_3_is_taken = _RAND_80[0:0];
  _RAND_81 = {1{`RANDOM}};
  rob_info_3_predict_miss = _RAND_81[0:0];
  _RAND_82 = {1{`RANDOM}};
  rob_info_3_gh_info = _RAND_82[3:0];
  _RAND_83 = {1{`RANDOM}};
  rob_info_3_op1_ready = _RAND_83[0:0];
  _RAND_84 = {1{`RANDOM}};
  rob_info_3_op1_tag = _RAND_84[2:0];
  _RAND_85 = {1{`RANDOM}};
  rob_info_3_op1_data = _RAND_85[31:0];
  _RAND_86 = {1{`RANDOM}};
  rob_info_3_op2_ready = _RAND_86[0:0];
  _RAND_87 = {1{`RANDOM}};
  rob_info_3_op2_tag = _RAND_87[2:0];
  _RAND_88 = {1{`RANDOM}};
  rob_info_3_op2_data = _RAND_88[31:0];
  _RAND_89 = {1{`RANDOM}};
  rob_info_3_imm_data = _RAND_89[31:0];
  _RAND_90 = {1{`RANDOM}};
  rob_info_3_is_init = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  rob_info_3_flush_on_commit = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  rob_info_4_is_valid = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  rob_info_4_busy = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  rob_info_4_uop = _RAND_94[5:0];
  _RAND_95 = {1{`RANDOM}};
  rob_info_4_unit_sel = _RAND_95[2:0];
  _RAND_96 = {1{`RANDOM}};
  rob_info_4_need_imm = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  rob_info_4_inst_addr = _RAND_97[31:0];
  _RAND_98 = {1{`RANDOM}};
  rob_info_4_commit_addr = _RAND_98[4:0];
  _RAND_99 = {1{`RANDOM}};
  rob_info_4_commit_data = _RAND_99[31:0];
  _RAND_100 = {1{`RANDOM}};
  rob_info_4_commit_ready = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  rob_info_4_is_branch = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  rob_info_4_predict_taken = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  rob_info_4_is_taken = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  rob_info_4_predict_miss = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  rob_info_4_gh_info = _RAND_105[3:0];
  _RAND_106 = {1{`RANDOM}};
  rob_info_4_op1_ready = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  rob_info_4_op1_tag = _RAND_107[2:0];
  _RAND_108 = {1{`RANDOM}};
  rob_info_4_op1_data = _RAND_108[31:0];
  _RAND_109 = {1{`RANDOM}};
  rob_info_4_op2_ready = _RAND_109[0:0];
  _RAND_110 = {1{`RANDOM}};
  rob_info_4_op2_tag = _RAND_110[2:0];
  _RAND_111 = {1{`RANDOM}};
  rob_info_4_op2_data = _RAND_111[31:0];
  _RAND_112 = {1{`RANDOM}};
  rob_info_4_imm_data = _RAND_112[31:0];
  _RAND_113 = {1{`RANDOM}};
  rob_info_4_is_init = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  rob_info_4_flush_on_commit = _RAND_114[0:0];
  _RAND_115 = {1{`RANDOM}};
  rob_info_5_is_valid = _RAND_115[0:0];
  _RAND_116 = {1{`RANDOM}};
  rob_info_5_busy = _RAND_116[0:0];
  _RAND_117 = {1{`RANDOM}};
  rob_info_5_uop = _RAND_117[5:0];
  _RAND_118 = {1{`RANDOM}};
  rob_info_5_unit_sel = _RAND_118[2:0];
  _RAND_119 = {1{`RANDOM}};
  rob_info_5_need_imm = _RAND_119[0:0];
  _RAND_120 = {1{`RANDOM}};
  rob_info_5_inst_addr = _RAND_120[31:0];
  _RAND_121 = {1{`RANDOM}};
  rob_info_5_commit_addr = _RAND_121[4:0];
  _RAND_122 = {1{`RANDOM}};
  rob_info_5_commit_data = _RAND_122[31:0];
  _RAND_123 = {1{`RANDOM}};
  rob_info_5_commit_ready = _RAND_123[0:0];
  _RAND_124 = {1{`RANDOM}};
  rob_info_5_is_branch = _RAND_124[0:0];
  _RAND_125 = {1{`RANDOM}};
  rob_info_5_predict_taken = _RAND_125[0:0];
  _RAND_126 = {1{`RANDOM}};
  rob_info_5_is_taken = _RAND_126[0:0];
  _RAND_127 = {1{`RANDOM}};
  rob_info_5_predict_miss = _RAND_127[0:0];
  _RAND_128 = {1{`RANDOM}};
  rob_info_5_gh_info = _RAND_128[3:0];
  _RAND_129 = {1{`RANDOM}};
  rob_info_5_op1_ready = _RAND_129[0:0];
  _RAND_130 = {1{`RANDOM}};
  rob_info_5_op1_tag = _RAND_130[2:0];
  _RAND_131 = {1{`RANDOM}};
  rob_info_5_op1_data = _RAND_131[31:0];
  _RAND_132 = {1{`RANDOM}};
  rob_info_5_op2_ready = _RAND_132[0:0];
  _RAND_133 = {1{`RANDOM}};
  rob_info_5_op2_tag = _RAND_133[2:0];
  _RAND_134 = {1{`RANDOM}};
  rob_info_5_op2_data = _RAND_134[31:0];
  _RAND_135 = {1{`RANDOM}};
  rob_info_5_imm_data = _RAND_135[31:0];
  _RAND_136 = {1{`RANDOM}};
  rob_info_5_is_init = _RAND_136[0:0];
  _RAND_137 = {1{`RANDOM}};
  rob_info_5_flush_on_commit = _RAND_137[0:0];
  _RAND_138 = {1{`RANDOM}};
  rob_info_6_is_valid = _RAND_138[0:0];
  _RAND_139 = {1{`RANDOM}};
  rob_info_6_busy = _RAND_139[0:0];
  _RAND_140 = {1{`RANDOM}};
  rob_info_6_uop = _RAND_140[5:0];
  _RAND_141 = {1{`RANDOM}};
  rob_info_6_unit_sel = _RAND_141[2:0];
  _RAND_142 = {1{`RANDOM}};
  rob_info_6_need_imm = _RAND_142[0:0];
  _RAND_143 = {1{`RANDOM}};
  rob_info_6_inst_addr = _RAND_143[31:0];
  _RAND_144 = {1{`RANDOM}};
  rob_info_6_commit_addr = _RAND_144[4:0];
  _RAND_145 = {1{`RANDOM}};
  rob_info_6_commit_data = _RAND_145[31:0];
  _RAND_146 = {1{`RANDOM}};
  rob_info_6_commit_ready = _RAND_146[0:0];
  _RAND_147 = {1{`RANDOM}};
  rob_info_6_is_branch = _RAND_147[0:0];
  _RAND_148 = {1{`RANDOM}};
  rob_info_6_predict_taken = _RAND_148[0:0];
  _RAND_149 = {1{`RANDOM}};
  rob_info_6_is_taken = _RAND_149[0:0];
  _RAND_150 = {1{`RANDOM}};
  rob_info_6_predict_miss = _RAND_150[0:0];
  _RAND_151 = {1{`RANDOM}};
  rob_info_6_gh_info = _RAND_151[3:0];
  _RAND_152 = {1{`RANDOM}};
  rob_info_6_op1_ready = _RAND_152[0:0];
  _RAND_153 = {1{`RANDOM}};
  rob_info_6_op1_tag = _RAND_153[2:0];
  _RAND_154 = {1{`RANDOM}};
  rob_info_6_op1_data = _RAND_154[31:0];
  _RAND_155 = {1{`RANDOM}};
  rob_info_6_op2_ready = _RAND_155[0:0];
  _RAND_156 = {1{`RANDOM}};
  rob_info_6_op2_tag = _RAND_156[2:0];
  _RAND_157 = {1{`RANDOM}};
  rob_info_6_op2_data = _RAND_157[31:0];
  _RAND_158 = {1{`RANDOM}};
  rob_info_6_imm_data = _RAND_158[31:0];
  _RAND_159 = {1{`RANDOM}};
  rob_info_6_is_init = _RAND_159[0:0];
  _RAND_160 = {1{`RANDOM}};
  rob_info_6_flush_on_commit = _RAND_160[0:0];
  _RAND_161 = {1{`RANDOM}};
  rob_info_7_is_valid = _RAND_161[0:0];
  _RAND_162 = {1{`RANDOM}};
  rob_info_7_busy = _RAND_162[0:0];
  _RAND_163 = {1{`RANDOM}};
  rob_info_7_uop = _RAND_163[5:0];
  _RAND_164 = {1{`RANDOM}};
  rob_info_7_unit_sel = _RAND_164[2:0];
  _RAND_165 = {1{`RANDOM}};
  rob_info_7_need_imm = _RAND_165[0:0];
  _RAND_166 = {1{`RANDOM}};
  rob_info_7_inst_addr = _RAND_166[31:0];
  _RAND_167 = {1{`RANDOM}};
  rob_info_7_commit_addr = _RAND_167[4:0];
  _RAND_168 = {1{`RANDOM}};
  rob_info_7_commit_data = _RAND_168[31:0];
  _RAND_169 = {1{`RANDOM}};
  rob_info_7_commit_ready = _RAND_169[0:0];
  _RAND_170 = {1{`RANDOM}};
  rob_info_7_is_branch = _RAND_170[0:0];
  _RAND_171 = {1{`RANDOM}};
  rob_info_7_predict_taken = _RAND_171[0:0];
  _RAND_172 = {1{`RANDOM}};
  rob_info_7_is_taken = _RAND_172[0:0];
  _RAND_173 = {1{`RANDOM}};
  rob_info_7_predict_miss = _RAND_173[0:0];
  _RAND_174 = {1{`RANDOM}};
  rob_info_7_gh_info = _RAND_174[3:0];
  _RAND_175 = {1{`RANDOM}};
  rob_info_7_op1_ready = _RAND_175[0:0];
  _RAND_176 = {1{`RANDOM}};
  rob_info_7_op1_tag = _RAND_176[2:0];
  _RAND_177 = {1{`RANDOM}};
  rob_info_7_op1_data = _RAND_177[31:0];
  _RAND_178 = {1{`RANDOM}};
  rob_info_7_op2_ready = _RAND_178[0:0];
  _RAND_179 = {1{`RANDOM}};
  rob_info_7_op2_tag = _RAND_179[2:0];
  _RAND_180 = {1{`RANDOM}};
  rob_info_7_op2_data = _RAND_180[31:0];
  _RAND_181 = {1{`RANDOM}};
  rob_info_7_imm_data = _RAND_181[31:0];
  _RAND_182 = {1{`RANDOM}};
  rob_info_7_is_init = _RAND_182[0:0];
  _RAND_183 = {1{`RANDOM}};
  rob_info_7_flush_on_commit = _RAND_183[0:0];
  _RAND_184 = {1{`RANDOM}};
  head = _RAND_184[7:0];
  _RAND_185 = {1{`RANDOM}};
  tail = _RAND_185[7:0];
  _RAND_186 = {1{`RANDOM}};
  maybe_full = _RAND_186[0:0];
  _RAND_187 = {1{`RANDOM}};
  waiting_delay = _RAND_187[0:0];
  _RAND_188 = {1{`RANDOM}};
  need_flush = _RAND_188[0:0];
  _RAND_189 = {1{`RANDOM}};
  rob_commit_1_des_rob = _RAND_189[2:0];
  _RAND_190 = {1{`RANDOM}};
  rob_commit_valid_1 = _RAND_190[0:0];
  _RAND_191 = {1{`RANDOM}};
  rob_commit_0_des_rob = _RAND_191[2:0];
  _RAND_192 = {1{`RANDOM}};
  rob_commit_valid_0 = _RAND_192[0:0];
  _RAND_193 = {1{`RANDOM}};
  rob_commit_1_commit_data = _RAND_193[31:0];
  _RAND_194 = {1{`RANDOM}};
  rob_commit_0_commit_data = _RAND_194[31:0];
  _RAND_195 = {1{`RANDOM}};
  rob_commit_0_commit_addr = _RAND_195[4:0];
  _RAND_196 = {1{`RANDOM}};
  rob_commit_1_commit_addr = _RAND_196[4:0];
  _RAND_197 = {1{`RANDOM}};
  branch_info_target_addr = _RAND_197[31:0];
  _RAND_198 = {1{`RANDOM}};
  branch_info_inst_addr = _RAND_198[31:0];
  _RAND_199 = {1{`RANDOM}};
  branch_info_gh_update = _RAND_199[3:0];
  _RAND_200 = {1{`RANDOM}};
  branch_info_is_branch = _RAND_200[0:0];
  _RAND_201 = {1{`RANDOM}};
  branch_info_is_taken = _RAND_201[0:0];
  _RAND_202 = {1{`RANDOM}};
  branch_info_predict_miss = _RAND_202[0:0];
  _RAND_203 = {1{`RANDOM}};
  branch_info_valid = _RAND_203[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Alu(
  input         clock,
  input         reset,
  input         io_dispatch_info_valid,
  input  [5:0]  io_dispatch_info_bits_uop,
  input         io_dispatch_info_bits_need_imm,
  input  [2:0]  io_dispatch_info_bits_rob_idx,
  input  [31:0] io_dispatch_info_bits_op1_data,
  input  [31:0] io_dispatch_info_bits_op2_data,
  input  [31:0] io_dispatch_info_bits_imm_data,
  output        io_wb_info_valid,
  output [2:0]  io_wb_info_bits_rob_idx,
  output [31:0] io_wb_info_bits_data,
  input         io_need_flush
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  reg [5:0] dispatch_info_uop; // @[Alu.scala 19:34]
  reg  dispatch_info_need_imm; // @[Alu.scala 19:34]
  reg [2:0] dispatch_info_rob_idx; // @[Alu.scala 19:34]
  reg [31:0] dispatch_info_op1_data; // @[Alu.scala 19:34]
  reg [31:0] dispatch_info_op2_data; // @[Alu.scala 19:34]
  reg [31:0] dispatch_info_imm_data; // @[Alu.scala 19:34]
  reg  dispatch_valid; // @[Alu.scala 21:38]
  wire [31:0] op2_data = dispatch_info_need_imm ? dispatch_info_imm_data : dispatch_info_op2_data; // @[Alu.scala 27:24]
  wire  _T_2 = 6'h1 == dispatch_info_uop; // @[Conditional.scala 37:30]
  wire [31:0] _result_data_T_1 = dispatch_info_op1_data + op2_data; // @[Alu.scala 33:31]
  wire  _T_5 = 6'h2 == dispatch_info_uop; // @[Conditional.scala 37:30]
  wire  _T_8 = 6'h3 == dispatch_info_uop; // @[Conditional.scala 37:30]
  wire [31:0] _result_data_T_5 = dispatch_info_op1_data - op2_data; // @[Alu.scala 39:31]
  wire  _T_11 = 6'h4 == dispatch_info_uop; // @[Conditional.scala 37:30]
  wire  _T_14 = 6'h5 == dispatch_info_uop; // @[Conditional.scala 37:30]
  wire [62:0] _GEN_42 = {{31'd0}, dispatch_info_op1_data}; // @[Alu.scala 45:40]
  wire [62:0] _result_data_T_9 = _GEN_42 << op2_data[4:0]; // @[Alu.scala 45:40]
  wire  _T_17 = 6'h6 == dispatch_info_uop; // @[Conditional.scala 37:30]
  wire [31:0] _result_data_T_11 = dispatch_info_op1_data >> op2_data[4:0]; // @[Alu.scala 48:41]
  wire  _T_20 = 6'h7 == dispatch_info_uop; // @[Conditional.scala 37:30]
  wire [31:0] _result_data_T_12 = dispatch_info_op1_data; // @[Alu.scala 51:38]
  wire [31:0] _result_data_T_14 = $signed(dispatch_info_op1_data) >>> op2_data; // @[Alu.scala 51:60]
  wire  _T_23 = 6'h8 == dispatch_info_uop; // @[Conditional.scala 37:30]
  wire [31:0] _result_data_T_16 = dispatch_info_need_imm ? dispatch_info_imm_data : dispatch_info_op2_data; // @[Alu.scala 54:58]
  wire  _T_26 = 6'h9 == dispatch_info_uop; // @[Conditional.scala 37:30]
  wire  _T_29 = 6'ha == dispatch_info_uop; // @[Conditional.scala 37:30]
  wire [31:0] _result_data_T_19 = dispatch_info_op1_data ^ op2_data; // @[Alu.scala 60:31]
  wire  _T_32 = 6'hb == dispatch_info_uop; // @[Conditional.scala 37:30]
  wire [31:0] _result_data_T_20 = dispatch_info_op1_data | op2_data; // @[Alu.scala 63:31]
  wire  _T_35 = 6'hc == dispatch_info_uop; // @[Conditional.scala 37:30]
  wire [31:0] _result_data_T_21 = dispatch_info_op1_data & op2_data; // @[Alu.scala 66:31]
  wire  _T_38 = 6'hd == dispatch_info_uop; // @[Conditional.scala 37:30]
  wire [15:0] result_data_hi = op2_data[15:0]; // @[Alu.scala 69:34]
  wire [31:0] _result_data_T_22 = {result_data_hi,16'h0}; // @[Cat.scala 30:58]
  wire  _T_41 = 6'he == dispatch_info_uop; // @[Conditional.scala 37:30]
  wire [31:0] _result_data_T_24 = ~_result_data_T_20; // @[Alu.scala 72:44]
  wire [31:0] _GEN_0 = _T_41 ? _result_data_T_24 : 32'h0; // @[Conditional.scala 39:67 Alu.scala 72:19 Alu.scala 30:15]
  wire [31:0] _GEN_1 = _T_38 ? _result_data_T_22 : _GEN_0; // @[Conditional.scala 39:67 Alu.scala 69:19]
  wire [31:0] _GEN_2 = _T_35 ? _result_data_T_21 : _GEN_1; // @[Conditional.scala 39:67 Alu.scala 66:19]
  wire [31:0] _GEN_3 = _T_32 ? _result_data_T_20 : _GEN_2; // @[Conditional.scala 39:67 Alu.scala 63:19]
  wire [31:0] _GEN_4 = _T_29 ? _result_data_T_19 : _GEN_3; // @[Conditional.scala 39:67 Alu.scala 60:19]
  wire [31:0] _GEN_5 = _T_26 ? {{31'd0}, dispatch_info_op1_data < op2_data} : _GEN_4; // @[Conditional.scala 39:67 Alu.scala 57:19]
  wire [31:0] _GEN_6 = _T_23 ? {{31'd0}, $signed(_result_data_T_12) < $signed(_result_data_T_16)} : _GEN_5; // @[Conditional.scala 39:67 Alu.scala 54:19]
  wire [31:0] _GEN_7 = _T_20 ? _result_data_T_14 : _GEN_6; // @[Conditional.scala 39:67 Alu.scala 51:19]
  wire [31:0] _GEN_8 = _T_17 ? _result_data_T_11 : _GEN_7; // @[Conditional.scala 39:67 Alu.scala 48:19]
  wire [62:0] _GEN_9 = _T_14 ? _result_data_T_9 : {{31'd0}, _GEN_8}; // @[Conditional.scala 39:67 Alu.scala 45:19]
  wire [62:0] _GEN_10 = _T_11 ? {{31'd0}, _result_data_T_5} : _GEN_9; // @[Conditional.scala 39:67 Alu.scala 42:19]
  wire [62:0] _GEN_11 = _T_8 ? {{31'd0}, _result_data_T_5} : _GEN_10; // @[Conditional.scala 39:67 Alu.scala 39:19]
  wire [62:0] _GEN_12 = _T_5 ? {{31'd0}, _result_data_T_1} : _GEN_11; // @[Conditional.scala 39:67 Alu.scala 36:19]
  wire [62:0] _GEN_13 = _T_2 ? {{31'd0}, _result_data_T_1} : _GEN_12; // @[Conditional.scala 40:58 Alu.scala 33:19]
  assign io_wb_info_valid = dispatch_valid; // @[Alu.scala 92:19]
  assign io_wb_info_bits_rob_idx = dispatch_info_rob_idx; // @[Alu.scala 88:26]
  assign io_wb_info_bits_data = _GEN_13[31:0]; // @[Alu.scala 28:25]
  always @(posedge clock) begin
    if (reset) begin // @[Alu.scala 102:23]
      dispatch_info_uop <= 6'h0; // @[Rob.scala 142:19]
    end else if (io_need_flush) begin // @[Alu.scala 95:22]
      dispatch_info_uop <= 6'h0; // @[Rob.scala 142:19]
    end else begin
      dispatch_info_uop <= io_dispatch_info_bits_uop; // @[Alu.scala 20:17]
    end
    if (reset) begin // @[Alu.scala 102:23]
      dispatch_info_need_imm <= 1'h0; // @[Rob.scala 143:19]
    end else if (io_need_flush) begin // @[Alu.scala 95:22]
      dispatch_info_need_imm <= 1'h0; // @[Rob.scala 143:19]
    end else begin
      dispatch_info_need_imm <= io_dispatch_info_bits_need_imm; // @[Alu.scala 20:17]
    end
    if (reset) begin // @[Alu.scala 102:23]
      dispatch_info_rob_idx <= 3'h0; // @[Rob.scala 144:19]
    end else if (io_need_flush) begin // @[Alu.scala 95:22]
      dispatch_info_rob_idx <= 3'h0; // @[Rob.scala 144:19]
    end else begin
      dispatch_info_rob_idx <= io_dispatch_info_bits_rob_idx; // @[Alu.scala 20:17]
    end
    if (reset) begin // @[Alu.scala 102:23]
      dispatch_info_op1_data <= 32'h0; // @[Rob.scala 146:19]
    end else if (io_need_flush) begin // @[Alu.scala 95:22]
      dispatch_info_op1_data <= 32'h0; // @[Rob.scala 146:19]
    end else begin
      dispatch_info_op1_data <= io_dispatch_info_bits_op1_data; // @[Alu.scala 20:17]
    end
    if (reset) begin // @[Alu.scala 102:23]
      dispatch_info_op2_data <= 32'h0; // @[Rob.scala 147:19]
    end else if (io_need_flush) begin // @[Alu.scala 95:22]
      dispatch_info_op2_data <= 32'h0; // @[Rob.scala 147:19]
    end else begin
      dispatch_info_op2_data <= io_dispatch_info_bits_op2_data; // @[Alu.scala 20:17]
    end
    if (reset) begin // @[Alu.scala 102:23]
      dispatch_info_imm_data <= 32'h0; // @[Rob.scala 148:19]
    end else if (io_need_flush) begin // @[Alu.scala 95:22]
      dispatch_info_imm_data <= 32'h0; // @[Rob.scala 148:19]
    end else begin
      dispatch_info_imm_data <= io_dispatch_info_bits_imm_data; // @[Alu.scala 20:17]
    end
    if (reset) begin // @[Alu.scala 21:38]
      dispatch_valid <= 1'h0; // @[Alu.scala 21:38]
    end else if (io_need_flush) begin // @[Alu.scala 95:22]
      dispatch_valid <= 1'h0; // @[Alu.scala 97:19]
    end else begin
      dispatch_valid <= io_dispatch_info_valid; // @[Alu.scala 22:17]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  dispatch_info_uop = _RAND_0[5:0];
  _RAND_1 = {1{`RANDOM}};
  dispatch_info_need_imm = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  dispatch_info_rob_idx = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  dispatch_info_op1_data = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  dispatch_info_op2_data = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  dispatch_info_imm_data = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  dispatch_valid = _RAND_6[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Bju(
  input         clock,
  input         reset,
  input         io_dispatch_info_valid,
  input  [5:0]  io_dispatch_info_bits_uop,
  input  [2:0]  io_dispatch_info_bits_rob_idx,
  input  [31:0] io_dispatch_info_bits_inst_addr,
  input  [31:0] io_dispatch_info_bits_op1_data,
  input  [31:0] io_dispatch_info_bits_op2_data,
  input  [31:0] io_dispatch_info_bits_imm_data,
  input         io_dispatch_info_bits_predict_taken,
  output        io_wb_info_valid,
  output [2:0]  io_wb_info_bits_rob_idx,
  output [31:0] io_wb_info_bits_data,
  output [31:0] io_wb_info_bits_target_addr,
  output        io_wb_info_bits_is_taken,
  output        io_wb_info_bits_predict_miss,
  input         io_need_flush
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg [5:0] dispatch_info_uop; // @[Bju.scala 21:34]
  reg [2:0] dispatch_info_rob_idx; // @[Bju.scala 21:34]
  reg [31:0] dispatch_info_inst_addr; // @[Bju.scala 21:34]
  reg [31:0] dispatch_info_op1_data; // @[Bju.scala 21:34]
  reg [31:0] dispatch_info_op2_data; // @[Bju.scala 21:34]
  reg [31:0] dispatch_info_imm_data; // @[Bju.scala 21:34]
  reg  dispatch_info_predict_taken; // @[Bju.scala 21:34]
  reg  dispatch_valid; // @[Bju.scala 23:38]
  wire [31:0] next_addr = dispatch_info_inst_addr + 32'h8; // @[Bju.scala 28:42]
  wire [29:0] branch_addr_hi = dispatch_info_imm_data[29:0]; // @[Bju.scala 29:81]
  wire [31:0] _branch_addr_T_2 = {branch_addr_hi,2'h0}; // @[Bju.scala 29:105]
  wire [31:0] _branch_addr_T_5 = $signed(dispatch_info_inst_addr) + $signed(_branch_addr_T_2); // @[Bju.scala 29:54]
  wire [31:0] branch_addr = $signed(_branch_addr_T_5) + 32'sh4; // @[Bju.scala 29:125]
  wire [3:0] jump_addr_hi_hi = dispatch_info_inst_addr[31:28]; // @[Bju.scala 30:46]
  wire [25:0] jump_addr_hi_lo = dispatch_info_imm_data[25:0]; // @[Bju.scala 30:76]
  wire [31:0] jump_addr = {jump_addr_hi_hi,jump_addr_hi_lo,2'h0}; // @[Cat.scala 30:58]
  wire  eq = dispatch_info_op1_data == dispatch_info_op2_data; // @[Bju.scala 33:32]
  wire  ez = dispatch_info_op1_data == 32'h0; // @[Bju.scala 34:34]
  wire  ltz = $signed(dispatch_info_op1_data) < 32'sh0; // @[Bju.scala 35:42]
  wire  _T_2 = 6'h18 == dispatch_info_uop; // @[Conditional.scala 37:30]
  wire  _T_5 = 6'h19 == dispatch_info_uop; // @[Conditional.scala 37:30]
  wire  _T_8 = 6'h1a == dispatch_info_uop; // @[Conditional.scala 37:30]
  wire  _T_11 = 6'h1b == dispatch_info_uop; // @[Conditional.scala 37:30]
  wire  _T_14 = 6'h1c == dispatch_info_uop; // @[Conditional.scala 37:30]
  wire  _T_17 = 6'h1d == dispatch_info_uop; // @[Conditional.scala 37:30]
  wire  _T_20 = 6'h1e == dispatch_info_uop; // @[Conditional.scala 37:30]
  wire  _T_23 = 6'h1f == dispatch_info_uop; // @[Conditional.scala 37:30]
  wire  _is_taken_T_2 = ~ltz; // @[Bju.scala 71:18]
  wire  _is_taken_T_4 = ~ltz & ~ez; // @[Bju.scala 71:23]
  wire  _T_26 = 6'h20 == dispatch_info_uop; // @[Conditional.scala 37:30]
  wire  _T_29 = 6'h21 == dispatch_info_uop; // @[Conditional.scala 37:30]
  wire  _T_32 = 6'h22 == dispatch_info_uop; // @[Conditional.scala 37:30]
  wire  _T_35 = 6'h23 == dispatch_info_uop; // @[Conditional.scala 37:30]
  wire  _GEN_0 = _T_35 & ltz; // @[Conditional.scala 39:67 Bju.scala 87:15 Bju.scala 39:11]
  wire [31:0] _GEN_1 = _T_35 ? branch_addr : 32'h0; // @[Conditional.scala 39:67 Bju.scala 88:18 Bju.scala 40:14]
  wire  _GEN_2 = _T_32 ? _is_taken_T_4 : _GEN_0; // @[Conditional.scala 39:67 Bju.scala 83:15]
  wire [31:0] _GEN_3 = _T_32 ? branch_addr : _GEN_1; // @[Conditional.scala 39:67 Bju.scala 84:18]
  wire  _GEN_4 = _T_29 ? _is_taken_T_2 : _GEN_2; // @[Conditional.scala 39:67 Bju.scala 79:15]
  wire [31:0] _GEN_5 = _T_29 ? branch_addr : _GEN_3; // @[Conditional.scala 39:67 Bju.scala 80:18]
  wire  _GEN_6 = _T_26 ? ltz : _GEN_4; // @[Conditional.scala 39:67 Bju.scala 75:15]
  wire [31:0] _GEN_7 = _T_26 ? branch_addr : _GEN_5; // @[Conditional.scala 39:67 Bju.scala 76:18]
  wire  _GEN_8 = _T_23 ? ~ltz & ~ez : _GEN_6; // @[Conditional.scala 39:67 Bju.scala 71:15]
  wire [31:0] _GEN_9 = _T_23 ? branch_addr : _GEN_7; // @[Conditional.scala 39:67 Bju.scala 72:18]
  wire  _GEN_10 = _T_20 ? ltz | ez : _GEN_8; // @[Conditional.scala 39:67 Bju.scala 67:15]
  wire [31:0] _GEN_11 = _T_20 ? branch_addr : _GEN_9; // @[Conditional.scala 39:67 Bju.scala 68:18]
  wire  _GEN_12 = _T_17 ? ~eq : _GEN_10; // @[Conditional.scala 39:67 Bju.scala 63:15]
  wire [31:0] _GEN_13 = _T_17 ? branch_addr : _GEN_11; // @[Conditional.scala 39:67 Bju.scala 64:18]
  wire  _GEN_14 = _T_14 ? eq : _GEN_12; // @[Conditional.scala 39:67 Bju.scala 59:15]
  wire [31:0] _GEN_15 = _T_14 ? branch_addr : _GEN_13; // @[Conditional.scala 39:67 Bju.scala 60:18]
  wire  _GEN_16 = _T_11 | _GEN_14; // @[Conditional.scala 39:67 Bju.scala 55:15]
  wire [31:0] _GEN_17 = _T_11 ? dispatch_info_op1_data : _GEN_15; // @[Conditional.scala 39:67 Bju.scala 56:18]
  wire  _GEN_18 = _T_8 | _GEN_16; // @[Conditional.scala 39:67 Bju.scala 51:15]
  wire [31:0] _GEN_19 = _T_8 ? dispatch_info_op1_data : _GEN_17; // @[Conditional.scala 39:67 Bju.scala 52:18]
  wire  _GEN_20 = _T_5 | _GEN_18; // @[Conditional.scala 39:67 Bju.scala 47:15]
  wire [31:0] _GEN_21 = _T_5 ? jump_addr : _GEN_19; // @[Conditional.scala 39:67 Bju.scala 48:18]
  wire  is_taken = _T_2 | _GEN_20; // @[Conditional.scala 40:58 Bju.scala 43:15]
  wire [31:0] target_addr = _T_2 ? jump_addr : _GEN_21; // @[Conditional.scala 40:58 Bju.scala 44:18]
  assign io_wb_info_valid = dispatch_valid; // @[Bju.scala 94:19]
  assign io_wb_info_bits_rob_idx = dispatch_info_rob_idx; // @[Bju.scala 97:26]
  assign io_wb_info_bits_data = dispatch_info_inst_addr + 32'h8; // @[Bju.scala 28:42]
  assign io_wb_info_bits_target_addr = ~is_taken & dispatch_info_predict_taken ? next_addr : target_addr; // @[Bju.scala 96:35]
  assign io_wb_info_bits_is_taken = _T_2 | _GEN_20; // @[Conditional.scala 40:58 Bju.scala 43:15]
  assign io_wb_info_bits_predict_miss = is_taken ^ dispatch_info_predict_taken; // @[Bju.scala 99:41]
  always @(posedge clock) begin
    if (reset) begin // @[Bju.scala 106:23]
      dispatch_info_uop <= 6'h0; // @[Rob.scala 142:19]
    end else if (io_need_flush) begin // @[Bju.scala 101:22]
      dispatch_info_uop <= 6'h0; // @[Rob.scala 142:19]
    end else begin
      dispatch_info_uop <= io_dispatch_info_bits_uop; // @[Bju.scala 22:17]
    end
    if (reset) begin // @[Bju.scala 106:23]
      dispatch_info_rob_idx <= 3'h0; // @[Rob.scala 144:19]
    end else if (io_need_flush) begin // @[Bju.scala 101:22]
      dispatch_info_rob_idx <= 3'h0; // @[Rob.scala 144:19]
    end else begin
      dispatch_info_rob_idx <= io_dispatch_info_bits_rob_idx; // @[Bju.scala 22:17]
    end
    if (reset) begin // @[Bju.scala 106:23]
      dispatch_info_inst_addr <= 32'h0; // @[Rob.scala 145:19]
    end else if (io_need_flush) begin // @[Bju.scala 101:22]
      dispatch_info_inst_addr <= 32'h0; // @[Rob.scala 145:19]
    end else begin
      dispatch_info_inst_addr <= io_dispatch_info_bits_inst_addr; // @[Bju.scala 22:17]
    end
    if (reset) begin // @[Bju.scala 106:23]
      dispatch_info_op1_data <= 32'h0; // @[Rob.scala 146:19]
    end else if (io_need_flush) begin // @[Bju.scala 101:22]
      dispatch_info_op1_data <= 32'h0; // @[Rob.scala 146:19]
    end else begin
      dispatch_info_op1_data <= io_dispatch_info_bits_op1_data; // @[Bju.scala 22:17]
    end
    if (reset) begin // @[Bju.scala 106:23]
      dispatch_info_op2_data <= 32'h0; // @[Rob.scala 147:19]
    end else if (io_need_flush) begin // @[Bju.scala 101:22]
      dispatch_info_op2_data <= 32'h0; // @[Rob.scala 147:19]
    end else begin
      dispatch_info_op2_data <= io_dispatch_info_bits_op2_data; // @[Bju.scala 22:17]
    end
    if (reset) begin // @[Bju.scala 106:23]
      dispatch_info_imm_data <= 32'h0; // @[Rob.scala 148:19]
    end else if (io_need_flush) begin // @[Bju.scala 101:22]
      dispatch_info_imm_data <= 32'h0; // @[Rob.scala 148:19]
    end else begin
      dispatch_info_imm_data <= io_dispatch_info_bits_imm_data; // @[Bju.scala 22:17]
    end
    if (reset) begin // @[Bju.scala 106:23]
      dispatch_info_predict_taken <= 1'h0; // @[Rob.scala 149:19]
    end else if (io_need_flush) begin // @[Bju.scala 101:22]
      dispatch_info_predict_taken <= 1'h0; // @[Rob.scala 149:19]
    end else begin
      dispatch_info_predict_taken <= io_dispatch_info_bits_predict_taken; // @[Bju.scala 22:17]
    end
    if (reset) begin // @[Bju.scala 23:38]
      dispatch_valid <= 1'h0; // @[Bju.scala 23:38]
    end else if (io_need_flush) begin // @[Bju.scala 101:22]
      dispatch_valid <= 1'h0; // @[Bju.scala 103:19]
    end else begin
      dispatch_valid <= io_dispatch_info_valid; // @[Bju.scala 24:17]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  dispatch_info_uop = _RAND_0[5:0];
  _RAND_1 = {1{`RANDOM}};
  dispatch_info_rob_idx = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  dispatch_info_inst_addr = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  dispatch_info_op1_data = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  dispatch_info_op2_data = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  dispatch_info_imm_data = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  dispatch_info_predict_taken = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  dispatch_valid = _RAND_7[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Lsu(
  input         clock,
  input         reset,
  output        io_dispatch_info_ready,
  input         io_dispatch_info_valid,
  input  [5:0]  io_dispatch_info_bits_uop,
  input  [2:0]  io_dispatch_info_bits_rob_idx,
  input  [31:0] io_dispatch_info_bits_op1_data,
  input  [31:0] io_dispatch_info_bits_op2_data,
  input  [31:0] io_dispatch_info_bits_imm_data,
  output        io_wb_info_valid,
  output [2:0]  io_wb_info_bits_rob_idx,
  output [31:0] io_wb_info_bits_data,
  input         io_rob_commit_0_valid,
  input  [2:0]  io_rob_commit_0_bits_des_rob,
  input         io_rob_commit_1_valid,
  input  [2:0]  io_rob_commit_1_bits_des_rob,
  input         io_cache_read_ready,
  output        io_cache_read_valid,
  output [31:0] io_cache_read_bits_addr,
  output [3:0]  io_cache_read_bits_rob_idx,
  input         io_cache_write_ready,
  output        io_cache_write_valid,
  output [31:0] io_cache_write_bits_addr,
  output [31:0] io_cache_write_bits_data,
  output [3:0]  io_cache_write_bits_byte_mask,
  input  [31:0] io_cache_resp_data,
  input         io_need_flush
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
`endif // RANDOMIZE_REG_INIT
  reg [5:0] dispatch_info_uop; // @[Lsu.scala 68:34]
  reg [2:0] dispatch_info_rob_idx; // @[Lsu.scala 68:34]
  reg [31:0] dispatch_info_op1_data; // @[Lsu.scala 68:34]
  reg [31:0] dispatch_info_op2_data; // @[Lsu.scala 68:34]
  reg [31:0] dispatch_info_imm_data; // @[Lsu.scala 68:34]
  reg  dispatch_valid; // @[Lsu.scala 69:38]
  reg [3:0] write_buffer_0_rob_idx; // @[Lsu.scala 70:34]
  reg [31:0] write_buffer_0_addr; // @[Lsu.scala 70:34]
  reg [31:0] write_buffer_0_data; // @[Lsu.scala 70:34]
  reg [3:0] write_buffer_0_byte_mask; // @[Lsu.scala 70:34]
  reg [3:0] write_buffer_1_rob_idx; // @[Lsu.scala 70:34]
  reg [31:0] write_buffer_1_addr; // @[Lsu.scala 70:34]
  reg [31:0] write_buffer_1_data; // @[Lsu.scala 70:34]
  reg [3:0] write_buffer_1_byte_mask; // @[Lsu.scala 70:34]
  reg [3:0] write_buffer_2_rob_idx; // @[Lsu.scala 70:34]
  reg [31:0] write_buffer_2_addr; // @[Lsu.scala 70:34]
  reg [31:0] write_buffer_2_data; // @[Lsu.scala 70:34]
  reg [3:0] write_buffer_2_byte_mask; // @[Lsu.scala 70:34]
  reg [3:0] write_buffer_3_rob_idx; // @[Lsu.scala 70:34]
  reg [31:0] write_buffer_3_addr; // @[Lsu.scala 70:34]
  reg [31:0] write_buffer_3_data; // @[Lsu.scala 70:34]
  reg [3:0] write_buffer_3_byte_mask; // @[Lsu.scala 70:34]
  reg  write_buffer_valid_0; // @[Lsu.scala 71:38]
  reg  write_buffer_valid_1; // @[Lsu.scala 71:38]
  reg  write_buffer_valid_2; // @[Lsu.scala 71:38]
  reg  write_buffer_valid_3; // @[Lsu.scala 71:38]
  reg  write_buffer_waiting_0; // @[Lsu.scala 72:38]
  reg  write_buffer_waiting_1; // @[Lsu.scala 72:38]
  reg  write_buffer_waiting_2; // @[Lsu.scala 72:38]
  reg  write_buffer_waiting_3; // @[Lsu.scala 72:38]
  reg  write_buffer_complete_0; // @[Lsu.scala 73:38]
  reg  write_buffer_complete_1; // @[Lsu.scala 73:38]
  reg  write_buffer_complete_2; // @[Lsu.scala 73:38]
  reg  write_buffer_complete_3; // @[Lsu.scala 73:38]
  reg  write_buffer_uncache_0; // @[Lsu.scala 74:38]
  reg  write_buffer_uncache_1; // @[Lsu.scala 74:38]
  reg  write_buffer_uncache_2; // @[Lsu.scala 74:38]
  reg  write_buffer_uncache_3; // @[Lsu.scala 74:38]
  reg [3:0] complete_head; // @[Lsu.scala 75:38]
  reg [3:0] tail; // @[Lsu.scala 76:38]
  reg  maybe_full; // @[Lsu.scala 77:38]
  wire  full = complete_head == tail & maybe_full; // @[Lsu.scala 78:54]
  wire [31:0] mem_addr = $signed(dispatch_info_imm_data) + $signed(dispatch_info_op1_data); // @[Lsu.scala 82:105]
  wire  is_ld = 6'h27 == dispatch_info_uop | (6'h29 == dispatch_info_uop | (6'h28 == dispatch_info_uop | (6'h2b ==
    dispatch_info_uop | 6'h2a == dispatch_info_uop))); // @[Mux.scala 80:57]
  wire  is_st = 6'h24 == dispatch_info_uop | (6'h25 == dispatch_info_uop | 6'h26 == dispatch_info_uop); // @[Mux.scala 80:57]
  wire [3:0] _byte_mask_T_10 = 6'h2a == dispatch_info_uop ? 4'h1 : 4'h0; // @[Mux.scala 80:57]
  wire [3:0] _byte_mask_T_12 = 6'h2b == dispatch_info_uop ? 4'h1 : _byte_mask_T_10; // @[Mux.scala 80:57]
  wire [3:0] _byte_mask_T_14 = 6'h28 == dispatch_info_uop ? 4'h3 : _byte_mask_T_12; // @[Mux.scala 80:57]
  wire [3:0] _byte_mask_T_16 = 6'h29 == dispatch_info_uop ? 4'h3 : _byte_mask_T_14; // @[Mux.scala 80:57]
  wire [3:0] _byte_mask_T_18 = 6'h27 == dispatch_info_uop ? 4'hf : _byte_mask_T_16; // @[Mux.scala 80:57]
  wire [3:0] _byte_mask_T_20 = 6'h26 == dispatch_info_uop ? 4'h1 : _byte_mask_T_18; // @[Mux.scala 80:57]
  wire [3:0] _byte_mask_T_22 = 6'h25 == dispatch_info_uop ? 4'h3 : _byte_mask_T_20; // @[Mux.scala 80:57]
  wire  is_uncache = mem_addr[31:4] == 28'hbfd003f; // @[Lsu.scala 114:47]
  wire  do_enq = ~full & is_st & dispatch_valid & ~io_need_flush; // @[Lsu.scala 118:46]
  wire [1:0] enq_idx_hi = tail[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] enq_idx_lo = tail[1:0]; // @[OneHot.scala 31:18]
  wire  enq_idx_hi_1 = |enq_idx_hi; // @[OneHot.scala 32:14]
  wire [1:0] _enq_idx_T = enq_idx_hi | enq_idx_lo; // @[OneHot.scala 32:28]
  wire  enq_idx_lo_1 = _enq_idx_T[1]; // @[CircuitMath.scala 30:8]
  wire [1:0] enq_idx = {enq_idx_hi_1,enq_idx_lo_1}; // @[Cat.scala 30:58]
  wire [3:0] _write_buffer_enq_idx_rob_idx = {{1'd0}, dispatch_info_rob_idx}; // @[Lsu.scala 121:35 Lsu.scala 121:35]
  wire  _GEN_368 = 2'h0 == enq_idx; // @[Lsu.scala 125:33 Lsu.scala 125:33 Lsu.scala 71:38]
  wire  _GEN_16 = 2'h0 == enq_idx | write_buffer_valid_0; // @[Lsu.scala 125:33 Lsu.scala 125:33 Lsu.scala 71:38]
  wire  _GEN_369 = 2'h1 == enq_idx; // @[Lsu.scala 125:33 Lsu.scala 125:33 Lsu.scala 71:38]
  wire  _GEN_17 = 2'h1 == enq_idx | write_buffer_valid_1; // @[Lsu.scala 125:33 Lsu.scala 125:33 Lsu.scala 71:38]
  wire  _GEN_370 = 2'h2 == enq_idx; // @[Lsu.scala 125:33 Lsu.scala 125:33 Lsu.scala 71:38]
  wire  _GEN_18 = 2'h2 == enq_idx | write_buffer_valid_2; // @[Lsu.scala 125:33 Lsu.scala 125:33 Lsu.scala 71:38]
  wire  _GEN_371 = 2'h3 == enq_idx; // @[Lsu.scala 125:33 Lsu.scala 125:33 Lsu.scala 71:38]
  wire  _GEN_19 = 2'h3 == enq_idx | write_buffer_valid_3; // @[Lsu.scala 125:33 Lsu.scala 125:33 Lsu.scala 71:38]
  wire  _GEN_20 = _GEN_368 | write_buffer_waiting_0; // @[Lsu.scala 126:35 Lsu.scala 126:35 Lsu.scala 72:38]
  wire  _GEN_21 = _GEN_369 | write_buffer_waiting_1; // @[Lsu.scala 126:35 Lsu.scala 126:35 Lsu.scala 72:38]
  wire  _GEN_22 = _GEN_370 | write_buffer_waiting_2; // @[Lsu.scala 126:35 Lsu.scala 126:35 Lsu.scala 72:38]
  wire  _GEN_23 = _GEN_371 | write_buffer_waiting_3; // @[Lsu.scala 126:35 Lsu.scala 126:35 Lsu.scala 72:38]
  wire  _GEN_24 = 2'h0 == enq_idx ? 1'h0 : write_buffer_complete_0; // @[Lsu.scala 127:36 Lsu.scala 127:36 Lsu.scala 73:38]
  wire  _GEN_25 = 2'h1 == enq_idx ? 1'h0 : write_buffer_complete_1; // @[Lsu.scala 127:36 Lsu.scala 127:36 Lsu.scala 73:38]
  wire  _GEN_26 = 2'h2 == enq_idx ? 1'h0 : write_buffer_complete_2; // @[Lsu.scala 127:36 Lsu.scala 127:36 Lsu.scala 73:38]
  wire  _GEN_27 = 2'h3 == enq_idx ? 1'h0 : write_buffer_complete_3; // @[Lsu.scala 127:36 Lsu.scala 127:36 Lsu.scala 73:38]
  wire [2:0] tail_hi = tail[2:0]; // @[Lsu.scala 60:12]
  wire  tail_lo = tail[3]; // @[Lsu.scala 60:29]
  wire [3:0] _tail_T = {tail_hi,tail_lo}; // @[Cat.scala 30:58]
  wire  _GEN_48 = do_enq ? _GEN_16 : write_buffer_valid_0; // @[Lsu.scala 120:16 Lsu.scala 71:38]
  wire  _GEN_49 = do_enq ? _GEN_17 : write_buffer_valid_1; // @[Lsu.scala 120:16 Lsu.scala 71:38]
  wire  _GEN_50 = do_enq ? _GEN_18 : write_buffer_valid_2; // @[Lsu.scala 120:16 Lsu.scala 71:38]
  wire  _GEN_51 = do_enq ? _GEN_19 : write_buffer_valid_3; // @[Lsu.scala 120:16 Lsu.scala 71:38]
  wire  _GEN_52 = do_enq ? _GEN_20 : write_buffer_waiting_0; // @[Lsu.scala 120:16 Lsu.scala 72:38]
  wire  _GEN_53 = do_enq ? _GEN_21 : write_buffer_waiting_1; // @[Lsu.scala 120:16 Lsu.scala 72:38]
  wire  _GEN_54 = do_enq ? _GEN_22 : write_buffer_waiting_2; // @[Lsu.scala 120:16 Lsu.scala 72:38]
  wire  _GEN_55 = do_enq ? _GEN_23 : write_buffer_waiting_3; // @[Lsu.scala 120:16 Lsu.scala 72:38]
  wire  _GEN_56 = do_enq ? _GEN_24 : write_buffer_complete_0; // @[Lsu.scala 120:16 Lsu.scala 73:38]
  wire  _GEN_57 = do_enq ? _GEN_25 : write_buffer_complete_1; // @[Lsu.scala 120:16 Lsu.scala 73:38]
  wire  _GEN_58 = do_enq ? _GEN_26 : write_buffer_complete_2; // @[Lsu.scala 120:16 Lsu.scala 73:38]
  wire  _GEN_59 = do_enq ? _GEN_27 : write_buffer_complete_3; // @[Lsu.scala 120:16 Lsu.scala 73:38]
  reg [3:0] ready_deq_idxs_0; // @[Lsu.scala 133:31]
  wire [2:0] ready_deq_idxs_hi = ready_deq_idxs_0[2:0]; // @[Lsu.scala 60:12]
  wire  ready_deq_idxs_lo = ready_deq_idxs_0[3]; // @[Lsu.scala 60:29]
  wire [3:0] ready_deq_idxs_1 = {ready_deq_idxs_hi,ready_deq_idxs_lo}; // @[Cat.scala 30:58]
  wire [1:0] ready_deq_idxs_hi_1 = ready_deq_idxs_0[1:0]; // @[Lsu.scala 60:12]
  wire [1:0] ready_deq_idxs_lo_1 = ready_deq_idxs_0[3:2]; // @[Lsu.scala 60:29]
  wire [3:0] ready_deq_idxs_2 = {ready_deq_idxs_hi_1,ready_deq_idxs_lo_1}; // @[Cat.scala 30:58]
  wire  ready_idx_hi_1 = |ready_deq_idxs_lo_1; // @[OneHot.scala 32:14]
  wire [1:0] _ready_idx_T = ready_deq_idxs_lo_1 | ready_deq_idxs_hi_1; // @[OneHot.scala 32:28]
  wire  ready_idx_lo_1 = _ready_idx_T[1]; // @[CircuitMath.scala 30:8]
  wire [1:0] ready_idx = {ready_idx_hi_1,ready_idx_lo_1}; // @[Cat.scala 30:58]
  wire  _GEN_66 = 2'h1 == ready_idx ? write_buffer_waiting_1 : write_buffer_waiting_0; // @[Lsu.scala 142:44 Lsu.scala 142:44]
  wire  _GEN_67 = 2'h2 == ready_idx ? write_buffer_waiting_2 : _GEN_66; // @[Lsu.scala 142:44 Lsu.scala 142:44]
  wire  _GEN_68 = 2'h3 == ready_idx ? write_buffer_waiting_3 : _GEN_67; // @[Lsu.scala 142:44 Lsu.scala 142:44]
  wire  _GEN_70 = 2'h1 == ready_idx ? write_buffer_valid_1 : write_buffer_valid_0; // @[Lsu.scala 142:44 Lsu.scala 142:44]
  wire  _GEN_71 = 2'h2 == ready_idx ? write_buffer_valid_2 : _GEN_70; // @[Lsu.scala 142:44 Lsu.scala 142:44]
  wire  _GEN_72 = 2'h3 == ready_idx ? write_buffer_valid_3 : _GEN_71; // @[Lsu.scala 142:44 Lsu.scala 142:44]
  wire [3:0] _GEN_74 = 2'h1 == ready_idx ? write_buffer_1_rob_idx : write_buffer_0_rob_idx; // @[Lsu.scala 142:135 Lsu.scala 142:135]
  wire [3:0] _GEN_75 = 2'h2 == ready_idx ? write_buffer_2_rob_idx : _GEN_74; // @[Lsu.scala 142:135 Lsu.scala 142:135]
  wire [3:0] _GEN_76 = 2'h3 == ready_idx ? write_buffer_3_rob_idx : _GEN_75; // @[Lsu.scala 142:135 Lsu.scala 142:135]
  wire [3:0] _GEN_376 = {{1'd0}, io_rob_commit_0_bits_des_rob}; // @[Lsu.scala 142:135]
  wire  _GEN_377 = 2'h0 == ready_idx; // @[Lsu.scala 143:42 Lsu.scala 143:42]
  wire  _GEN_77 = 2'h0 == ready_idx | _GEN_56; // @[Lsu.scala 143:42 Lsu.scala 143:42]
  wire  _GEN_378 = 2'h1 == ready_idx; // @[Lsu.scala 143:42 Lsu.scala 143:42]
  wire  _GEN_78 = 2'h1 == ready_idx | _GEN_57; // @[Lsu.scala 143:42 Lsu.scala 143:42]
  wire  _GEN_379 = 2'h2 == ready_idx; // @[Lsu.scala 143:42 Lsu.scala 143:42]
  wire  _GEN_79 = 2'h2 == ready_idx | _GEN_58; // @[Lsu.scala 143:42 Lsu.scala 143:42]
  wire  _GEN_380 = 2'h3 == ready_idx; // @[Lsu.scala 143:42 Lsu.scala 143:42]
  wire  _GEN_80 = 2'h3 == ready_idx | _GEN_59; // @[Lsu.scala 143:42 Lsu.scala 143:42]
  wire  _GEN_81 = 2'h0 == ready_idx ? 1'h0 : _GEN_52; // @[Lsu.scala 144:41 Lsu.scala 144:41]
  wire  _GEN_82 = 2'h1 == ready_idx ? 1'h0 : _GEN_53; // @[Lsu.scala 144:41 Lsu.scala 144:41]
  wire  _GEN_83 = 2'h2 == ready_idx ? 1'h0 : _GEN_54; // @[Lsu.scala 144:41 Lsu.scala 144:41]
  wire  _GEN_84 = 2'h3 == ready_idx ? 1'h0 : _GEN_55; // @[Lsu.scala 144:41 Lsu.scala 144:41]
  wire  _GEN_89 = _GEN_68 & _GEN_72 & io_rob_commit_0_valid & _GEN_376 == _GEN_76 ? _GEN_77 : _GEN_56; // @[Lsu.scala 142:172]
  wire  _GEN_90 = _GEN_68 & _GEN_72 & io_rob_commit_0_valid & _GEN_376 == _GEN_76 ? _GEN_78 : _GEN_57; // @[Lsu.scala 142:172]
  wire  _GEN_91 = _GEN_68 & _GEN_72 & io_rob_commit_0_valid & _GEN_376 == _GEN_76 ? _GEN_79 : _GEN_58; // @[Lsu.scala 142:172]
  wire  _GEN_92 = _GEN_68 & _GEN_72 & io_rob_commit_0_valid & _GEN_376 == _GEN_76 ? _GEN_80 : _GEN_59; // @[Lsu.scala 142:172]
  wire  _GEN_93 = _GEN_68 & _GEN_72 & io_rob_commit_0_valid & _GEN_376 == _GEN_76 ? _GEN_81 : _GEN_52; // @[Lsu.scala 142:172]
  wire  _GEN_94 = _GEN_68 & _GEN_72 & io_rob_commit_0_valid & _GEN_376 == _GEN_76 ? _GEN_82 : _GEN_53; // @[Lsu.scala 142:172]
  wire  _GEN_95 = _GEN_68 & _GEN_72 & io_rob_commit_0_valid & _GEN_376 == _GEN_76 ? _GEN_83 : _GEN_54; // @[Lsu.scala 142:172]
  wire  _GEN_96 = _GEN_68 & _GEN_72 & io_rob_commit_0_valid & _GEN_376 == _GEN_76 ? _GEN_84 : _GEN_55; // @[Lsu.scala 142:172]
  wire  _GEN_98 = _GEN_68 & _GEN_72 & io_rob_commit_0_valid & _GEN_376 == _GEN_76 & _GEN_377; // @[Lsu.scala 142:172 Lsu.scala 136:30]
  wire  _GEN_99 = _GEN_68 & _GEN_72 & io_rob_commit_0_valid & _GEN_376 == _GEN_76 & _GEN_378; // @[Lsu.scala 142:172 Lsu.scala 136:30]
  wire  _GEN_100 = _GEN_68 & _GEN_72 & io_rob_commit_0_valid & _GEN_376 == _GEN_76 & _GEN_379; // @[Lsu.scala 142:172 Lsu.scala 136:30]
  wire  _GEN_101 = _GEN_68 & _GEN_72 & io_rob_commit_0_valid & _GEN_376 == _GEN_76 & _GEN_380; // @[Lsu.scala 142:172 Lsu.scala 136:30]
  wire [3:0] _GEN_381 = {{1'd0}, io_rob_commit_1_bits_des_rob}; // @[Lsu.scala 142:135]
  wire  _GEN_102 = 2'h0 == ready_idx | _GEN_89; // @[Lsu.scala 143:42 Lsu.scala 143:42]
  wire  _GEN_103 = 2'h1 == ready_idx | _GEN_90; // @[Lsu.scala 143:42 Lsu.scala 143:42]
  wire  _GEN_104 = 2'h2 == ready_idx | _GEN_91; // @[Lsu.scala 143:42 Lsu.scala 143:42]
  wire  _GEN_105 = 2'h3 == ready_idx | _GEN_92; // @[Lsu.scala 143:42 Lsu.scala 143:42]
  wire  _GEN_106 = 2'h0 == ready_idx ? 1'h0 : _GEN_93; // @[Lsu.scala 144:41 Lsu.scala 144:41]
  wire  _GEN_107 = 2'h1 == ready_idx ? 1'h0 : _GEN_94; // @[Lsu.scala 144:41 Lsu.scala 144:41]
  wire  _GEN_108 = 2'h2 == ready_idx ? 1'h0 : _GEN_95; // @[Lsu.scala 144:41 Lsu.scala 144:41]
  wire  _GEN_109 = 2'h3 == ready_idx ? 1'h0 : _GEN_96; // @[Lsu.scala 144:41 Lsu.scala 144:41]
  wire  _GEN_110 = _GEN_377 | _GEN_98; // @[Lsu.scala 146:33 Lsu.scala 146:33]
  wire  _GEN_111 = _GEN_378 | _GEN_99; // @[Lsu.scala 146:33 Lsu.scala 146:33]
  wire  _GEN_112 = _GEN_379 | _GEN_100; // @[Lsu.scala 146:33 Lsu.scala 146:33]
  wire  _GEN_113 = _GEN_380 | _GEN_101; // @[Lsu.scala 146:33 Lsu.scala 146:33]
  wire  _GEN_114 = _GEN_68 & _GEN_72 & io_rob_commit_1_valid & _GEN_381 == _GEN_76 ? _GEN_102 : _GEN_89; // @[Lsu.scala 142:172]
  wire  _GEN_115 = _GEN_68 & _GEN_72 & io_rob_commit_1_valid & _GEN_381 == _GEN_76 ? _GEN_103 : _GEN_90; // @[Lsu.scala 142:172]
  wire  _GEN_116 = _GEN_68 & _GEN_72 & io_rob_commit_1_valid & _GEN_381 == _GEN_76 ? _GEN_104 : _GEN_91; // @[Lsu.scala 142:172]
  wire  _GEN_117 = _GEN_68 & _GEN_72 & io_rob_commit_1_valid & _GEN_381 == _GEN_76 ? _GEN_105 : _GEN_92; // @[Lsu.scala 142:172]
  wire  _GEN_118 = _GEN_68 & _GEN_72 & io_rob_commit_1_valid & _GEN_381 == _GEN_76 ? _GEN_106 : _GEN_93; // @[Lsu.scala 142:172]
  wire  _GEN_119 = _GEN_68 & _GEN_72 & io_rob_commit_1_valid & _GEN_381 == _GEN_76 ? _GEN_107 : _GEN_94; // @[Lsu.scala 142:172]
  wire  _GEN_120 = _GEN_68 & _GEN_72 & io_rob_commit_1_valid & _GEN_381 == _GEN_76 ? _GEN_108 : _GEN_95; // @[Lsu.scala 142:172]
  wire  _GEN_121 = _GEN_68 & _GEN_72 & io_rob_commit_1_valid & _GEN_381 == _GEN_76 ? _GEN_109 : _GEN_96; // @[Lsu.scala 142:172]
  wire  ready_valid_0 = _GEN_68 & _GEN_72 & io_rob_commit_1_valid & _GEN_381 == _GEN_76 | _GEN_68 & _GEN_72 &
    io_rob_commit_0_valid & _GEN_376 == _GEN_76; // @[Lsu.scala 142:172 Lsu.scala 145:24]
  wire  _GEN_123 = _GEN_68 & _GEN_72 & io_rob_commit_1_valid & _GEN_381 == _GEN_76 ? _GEN_110 : _GEN_98; // @[Lsu.scala 142:172]
  wire  _GEN_124 = _GEN_68 & _GEN_72 & io_rob_commit_1_valid & _GEN_381 == _GEN_76 ? _GEN_111 : _GEN_99; // @[Lsu.scala 142:172]
  wire  _GEN_125 = _GEN_68 & _GEN_72 & io_rob_commit_1_valid & _GEN_381 == _GEN_76 ? _GEN_112 : _GEN_100; // @[Lsu.scala 142:172]
  wire  _GEN_126 = _GEN_68 & _GEN_72 & io_rob_commit_1_valid & _GEN_381 == _GEN_76 ? _GEN_113 : _GEN_101; // @[Lsu.scala 142:172]
  wire [1:0] ready_idx_hi_2 = ready_deq_idxs_1[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] ready_idx_lo_2 = ready_deq_idxs_1[1:0]; // @[OneHot.scala 31:18]
  wire  ready_idx_hi_3 = |ready_idx_hi_2; // @[OneHot.scala 32:14]
  wire [1:0] _ready_idx_T_1 = ready_idx_hi_2 | ready_idx_lo_2; // @[OneHot.scala 32:28]
  wire  ready_idx_lo_3 = _ready_idx_T_1[1]; // @[CircuitMath.scala 30:8]
  wire [1:0] ready_idx_1 = {ready_idx_hi_3,ready_idx_lo_3}; // @[Cat.scala 30:58]
  wire  _GEN_128 = 2'h1 == ready_idx_1 ? write_buffer_waiting_1 : write_buffer_waiting_0; // @[Lsu.scala 142:44 Lsu.scala 142:44]
  wire  _GEN_129 = 2'h2 == ready_idx_1 ? write_buffer_waiting_2 : _GEN_128; // @[Lsu.scala 142:44 Lsu.scala 142:44]
  wire  _GEN_130 = 2'h3 == ready_idx_1 ? write_buffer_waiting_3 : _GEN_129; // @[Lsu.scala 142:44 Lsu.scala 142:44]
  wire  _GEN_132 = 2'h1 == ready_idx_1 ? write_buffer_valid_1 : write_buffer_valid_0; // @[Lsu.scala 142:44 Lsu.scala 142:44]
  wire  _GEN_133 = 2'h2 == ready_idx_1 ? write_buffer_valid_2 : _GEN_132; // @[Lsu.scala 142:44 Lsu.scala 142:44]
  wire  _GEN_134 = 2'h3 == ready_idx_1 ? write_buffer_valid_3 : _GEN_133; // @[Lsu.scala 142:44 Lsu.scala 142:44]
  wire [3:0] _GEN_136 = 2'h1 == ready_idx_1 ? write_buffer_1_rob_idx : write_buffer_0_rob_idx; // @[Lsu.scala 142:135 Lsu.scala 142:135]
  wire [3:0] _GEN_137 = 2'h2 == ready_idx_1 ? write_buffer_2_rob_idx : _GEN_136; // @[Lsu.scala 142:135 Lsu.scala 142:135]
  wire [3:0] _GEN_138 = 2'h3 == ready_idx_1 ? write_buffer_3_rob_idx : _GEN_137; // @[Lsu.scala 142:135 Lsu.scala 142:135]
  wire  _GEN_391 = 2'h0 == ready_idx_1; // @[Lsu.scala 143:42 Lsu.scala 143:42]
  wire  _GEN_139 = 2'h0 == ready_idx_1 | _GEN_114; // @[Lsu.scala 143:42 Lsu.scala 143:42]
  wire  _GEN_392 = 2'h1 == ready_idx_1; // @[Lsu.scala 143:42 Lsu.scala 143:42]
  wire  _GEN_140 = 2'h1 == ready_idx_1 | _GEN_115; // @[Lsu.scala 143:42 Lsu.scala 143:42]
  wire  _GEN_393 = 2'h2 == ready_idx_1; // @[Lsu.scala 143:42 Lsu.scala 143:42]
  wire  _GEN_141 = 2'h2 == ready_idx_1 | _GEN_116; // @[Lsu.scala 143:42 Lsu.scala 143:42]
  wire  _GEN_394 = 2'h3 == ready_idx_1; // @[Lsu.scala 143:42 Lsu.scala 143:42]
  wire  _GEN_142 = 2'h3 == ready_idx_1 | _GEN_117; // @[Lsu.scala 143:42 Lsu.scala 143:42]
  wire  _GEN_143 = 2'h0 == ready_idx_1 ? 1'h0 : _GEN_118; // @[Lsu.scala 144:41 Lsu.scala 144:41]
  wire  _GEN_144 = 2'h1 == ready_idx_1 ? 1'h0 : _GEN_119; // @[Lsu.scala 144:41 Lsu.scala 144:41]
  wire  _GEN_145 = 2'h2 == ready_idx_1 ? 1'h0 : _GEN_120; // @[Lsu.scala 144:41 Lsu.scala 144:41]
  wire  _GEN_146 = 2'h3 == ready_idx_1 ? 1'h0 : _GEN_121; // @[Lsu.scala 144:41 Lsu.scala 144:41]
  wire  _GEN_147 = _GEN_391 | _GEN_123; // @[Lsu.scala 146:33 Lsu.scala 146:33]
  wire  _GEN_148 = _GEN_392 | _GEN_124; // @[Lsu.scala 146:33 Lsu.scala 146:33]
  wire  _GEN_149 = _GEN_393 | _GEN_125; // @[Lsu.scala 146:33 Lsu.scala 146:33]
  wire  _GEN_150 = _GEN_394 | _GEN_126; // @[Lsu.scala 146:33 Lsu.scala 146:33]
  wire  _GEN_151 = _GEN_130 & _GEN_134 & io_rob_commit_0_valid & _GEN_376 == _GEN_138 ? _GEN_139 : _GEN_114; // @[Lsu.scala 142:172]
  wire  _GEN_152 = _GEN_130 & _GEN_134 & io_rob_commit_0_valid & _GEN_376 == _GEN_138 ? _GEN_140 : _GEN_115; // @[Lsu.scala 142:172]
  wire  _GEN_153 = _GEN_130 & _GEN_134 & io_rob_commit_0_valid & _GEN_376 == _GEN_138 ? _GEN_141 : _GEN_116; // @[Lsu.scala 142:172]
  wire  _GEN_154 = _GEN_130 & _GEN_134 & io_rob_commit_0_valid & _GEN_376 == _GEN_138 ? _GEN_142 : _GEN_117; // @[Lsu.scala 142:172]
  wire  _GEN_155 = _GEN_130 & _GEN_134 & io_rob_commit_0_valid & _GEN_376 == _GEN_138 ? _GEN_143 : _GEN_118; // @[Lsu.scala 142:172]
  wire  _GEN_156 = _GEN_130 & _GEN_134 & io_rob_commit_0_valid & _GEN_376 == _GEN_138 ? _GEN_144 : _GEN_119; // @[Lsu.scala 142:172]
  wire  _GEN_157 = _GEN_130 & _GEN_134 & io_rob_commit_0_valid & _GEN_376 == _GEN_138 ? _GEN_145 : _GEN_120; // @[Lsu.scala 142:172]
  wire  _GEN_158 = _GEN_130 & _GEN_134 & io_rob_commit_0_valid & _GEN_376 == _GEN_138 ? _GEN_146 : _GEN_121; // @[Lsu.scala 142:172]
  wire  _GEN_160 = _GEN_130 & _GEN_134 & io_rob_commit_0_valid & _GEN_376 == _GEN_138 ? _GEN_147 : _GEN_123; // @[Lsu.scala 142:172]
  wire  _GEN_161 = _GEN_130 & _GEN_134 & io_rob_commit_0_valid & _GEN_376 == _GEN_138 ? _GEN_148 : _GEN_124; // @[Lsu.scala 142:172]
  wire  _GEN_162 = _GEN_130 & _GEN_134 & io_rob_commit_0_valid & _GEN_376 == _GEN_138 ? _GEN_149 : _GEN_125; // @[Lsu.scala 142:172]
  wire  _GEN_163 = _GEN_130 & _GEN_134 & io_rob_commit_0_valid & _GEN_376 == _GEN_138 ? _GEN_150 : _GEN_126; // @[Lsu.scala 142:172]
  wire  _GEN_164 = 2'h0 == ready_idx_1 | _GEN_151; // @[Lsu.scala 143:42 Lsu.scala 143:42]
  wire  _GEN_165 = 2'h1 == ready_idx_1 | _GEN_152; // @[Lsu.scala 143:42 Lsu.scala 143:42]
  wire  _GEN_166 = 2'h2 == ready_idx_1 | _GEN_153; // @[Lsu.scala 143:42 Lsu.scala 143:42]
  wire  _GEN_167 = 2'h3 == ready_idx_1 | _GEN_154; // @[Lsu.scala 143:42 Lsu.scala 143:42]
  wire  _GEN_168 = 2'h0 == ready_idx_1 ? 1'h0 : _GEN_155; // @[Lsu.scala 144:41 Lsu.scala 144:41]
  wire  _GEN_169 = 2'h1 == ready_idx_1 ? 1'h0 : _GEN_156; // @[Lsu.scala 144:41 Lsu.scala 144:41]
  wire  _GEN_170 = 2'h2 == ready_idx_1 ? 1'h0 : _GEN_157; // @[Lsu.scala 144:41 Lsu.scala 144:41]
  wire  _GEN_171 = 2'h3 == ready_idx_1 ? 1'h0 : _GEN_158; // @[Lsu.scala 144:41 Lsu.scala 144:41]
  wire  _GEN_172 = _GEN_391 | _GEN_160; // @[Lsu.scala 146:33 Lsu.scala 146:33]
  wire  _GEN_173 = _GEN_392 | _GEN_161; // @[Lsu.scala 146:33 Lsu.scala 146:33]
  wire  _GEN_174 = _GEN_393 | _GEN_162; // @[Lsu.scala 146:33 Lsu.scala 146:33]
  wire  _GEN_175 = _GEN_394 | _GEN_163; // @[Lsu.scala 146:33 Lsu.scala 146:33]
  wire  _GEN_180 = _GEN_130 & _GEN_134 & io_rob_commit_1_valid & _GEN_381 == _GEN_138 ? _GEN_168 : _GEN_155; // @[Lsu.scala 142:172]
  wire  _GEN_181 = _GEN_130 & _GEN_134 & io_rob_commit_1_valid & _GEN_381 == _GEN_138 ? _GEN_169 : _GEN_156; // @[Lsu.scala 142:172]
  wire  _GEN_182 = _GEN_130 & _GEN_134 & io_rob_commit_1_valid & _GEN_381 == _GEN_138 ? _GEN_170 : _GEN_157; // @[Lsu.scala 142:172]
  wire  _GEN_183 = _GEN_130 & _GEN_134 & io_rob_commit_1_valid & _GEN_381 == _GEN_138 ? _GEN_171 : _GEN_158; // @[Lsu.scala 142:172]
  wire  ready_valid_1 = _GEN_130 & _GEN_134 & io_rob_commit_1_valid & _GEN_381 == _GEN_138 | _GEN_130 & _GEN_134 &
    io_rob_commit_0_valid & _GEN_376 == _GEN_138; // @[Lsu.scala 142:172 Lsu.scala 145:24]
  wire  will_complete_0 = _GEN_130 & _GEN_134 & io_rob_commit_1_valid & _GEN_381 == _GEN_138 ? _GEN_172 : _GEN_160; // @[Lsu.scala 142:172]
  wire  will_complete_1 = _GEN_130 & _GEN_134 & io_rob_commit_1_valid & _GEN_381 == _GEN_138 ? _GEN_173 : _GEN_161; // @[Lsu.scala 142:172]
  wire  will_complete_2 = _GEN_130 & _GEN_134 & io_rob_commit_1_valid & _GEN_381 == _GEN_138 ? _GEN_174 : _GEN_162; // @[Lsu.scala 142:172]
  wire  will_complete_3 = _GEN_130 & _GEN_134 & io_rob_commit_1_valid & _GEN_381 == _GEN_138 ? _GEN_175 : _GEN_163; // @[Lsu.scala 142:172]
  wire [3:0] _T_18 = ready_valid_0 & ready_deq_idxs_0 != tail ? ready_deq_idxs_1 : ready_deq_idxs_0; // @[Lsu.scala 152:26]
  wire [1:0] complete_head_idx_hi = complete_head[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] complete_head_idx_lo = complete_head[1:0]; // @[OneHot.scala 31:18]
  wire  complete_head_idx_hi_1 = |complete_head_idx_hi; // @[OneHot.scala 32:14]
  wire [1:0] _complete_head_idx_T = complete_head_idx_hi | complete_head_idx_lo; // @[OneHot.scala 32:28]
  wire  complete_head_idx_lo_1 = _complete_head_idx_T[1]; // @[CircuitMath.scala 30:8]
  wire [1:0] complete_head_idx = {complete_head_idx_hi_1,complete_head_idx_lo_1}; // @[Cat.scala 30:58]
  wire  _GEN_190 = 2'h1 == complete_head_idx ? write_buffer_valid_1 : write_buffer_valid_0; // @[Lsu.scala 163:47 Lsu.scala 163:47]
  wire  _GEN_191 = 2'h2 == complete_head_idx ? write_buffer_valid_2 : _GEN_190; // @[Lsu.scala 163:47 Lsu.scala 163:47]
  wire  _GEN_192 = 2'h3 == complete_head_idx ? write_buffer_valid_3 : _GEN_191; // @[Lsu.scala 163:47 Lsu.scala 163:47]
  wire  _GEN_194 = 2'h1 == complete_head_idx ? write_buffer_complete_1 : write_buffer_complete_0; // @[Lsu.scala 163:47 Lsu.scala 163:47]
  wire  _GEN_195 = 2'h2 == complete_head_idx ? write_buffer_complete_2 : _GEN_194; // @[Lsu.scala 163:47 Lsu.scala 163:47]
  wire  _GEN_196 = 2'h3 == complete_head_idx ? write_buffer_complete_3 : _GEN_195; // @[Lsu.scala 163:47 Lsu.scala 163:47]
  wire [31:0] _GEN_198 = 2'h1 == complete_head_idx ? write_buffer_1_data : write_buffer_0_data; // @[Lsu.scala 164:28 Lsu.scala 164:28]
  wire [31:0] _GEN_199 = 2'h2 == complete_head_idx ? write_buffer_2_data : _GEN_198; // @[Lsu.scala 164:28 Lsu.scala 164:28]
  wire [31:0] _GEN_202 = 2'h1 == complete_head_idx ? write_buffer_1_addr : write_buffer_0_addr; // @[Lsu.scala 165:28 Lsu.scala 165:28]
  wire [31:0] _GEN_203 = 2'h2 == complete_head_idx ? write_buffer_2_addr : _GEN_202; // @[Lsu.scala 165:28 Lsu.scala 165:28]
  wire [3:0] _GEN_206 = 2'h1 == complete_head_idx ? write_buffer_1_byte_mask : write_buffer_0_byte_mask; // @[Lsu.scala 166:33 Lsu.scala 166:33]
  wire [3:0] _GEN_207 = 2'h2 == complete_head_idx ? write_buffer_2_byte_mask : _GEN_206; // @[Lsu.scala 166:33 Lsu.scala 166:33]
  wire [2:0] complete_head_hi = complete_head[2:0]; // @[Lsu.scala 60:12]
  wire  complete_head_lo = complete_head[3]; // @[Lsu.scala 60:29]
  wire [3:0] _complete_head_T = {complete_head_hi,complete_head_lo}; // @[Cat.scala 30:58]
  wire  _GEN_209 = 2'h0 == complete_head_idx ? 1'h0 : _GEN_48; // @[Lsu.scala 170:43 Lsu.scala 170:43]
  wire  _GEN_210 = 2'h1 == complete_head_idx ? 1'h0 : _GEN_49; // @[Lsu.scala 170:43 Lsu.scala 170:43]
  wire  _GEN_211 = 2'h2 == complete_head_idx ? 1'h0 : _GEN_50; // @[Lsu.scala 170:43 Lsu.scala 170:43]
  wire  _GEN_212 = 2'h3 == complete_head_idx ? 1'h0 : _GEN_51; // @[Lsu.scala 170:43 Lsu.scala 170:43]
  wire  _GEN_214 = io_cache_write_ready ? _GEN_209 : _GEN_48; // @[Lsu.scala 168:16]
  wire  _GEN_215 = io_cache_write_ready ? _GEN_210 : _GEN_49; // @[Lsu.scala 168:16]
  wire  _GEN_216 = io_cache_write_ready ? _GEN_211 : _GEN_50; // @[Lsu.scala 168:16]
  wire  _GEN_217 = io_cache_write_ready ? _GEN_212 : _GEN_51; // @[Lsu.scala 168:16]
  wire  _GEN_218 = io_cache_write_ready ? 1'h0 : maybe_full; // @[Lsu.scala 175:22 Lsu.scala 176:16 Lsu.scala 77:38]
  wire  _GEN_219 = do_enq | _GEN_218; // @[Lsu.scala 173:16 Lsu.scala 174:16]
  wire  do_read = dispatch_valid & is_ld; // @[Lsu.scala 179:40]
  wire [1:0] bypass_idxs_hi_3 = _tail_T[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] bypass_idxs_lo_3 = _tail_T[1:0]; // @[OneHot.scala 31:18]
  wire  bypass_idxs_hi_4 = |bypass_idxs_hi_3; // @[OneHot.scala 32:14]
  wire [1:0] _bypass_idxs_T_3 = bypass_idxs_hi_3 | bypass_idxs_lo_3; // @[OneHot.scala 32:28]
  wire  bypass_idxs_lo_4 = _bypass_idxs_T_3[1]; // @[CircuitMath.scala 30:8]
  wire [1:0] bypass_idxs_2 = {bypass_idxs_hi_4,bypass_idxs_lo_4}; // @[Cat.scala 30:58]
  wire [3:0] _bypass_idxs_T_5 = {enq_idx_lo,enq_idx_hi}; // @[Cat.scala 30:58]
  wire [1:0] bypass_idxs_hi_6 = _bypass_idxs_T_5[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] bypass_idxs_lo_6 = _bypass_idxs_T_5[1:0]; // @[OneHot.scala 31:18]
  wire  bypass_idxs_hi_7 = |bypass_idxs_hi_6; // @[OneHot.scala 32:14]
  wire [1:0] _bypass_idxs_T_6 = bypass_idxs_hi_6 | bypass_idxs_lo_6; // @[OneHot.scala 32:28]
  wire  bypass_idxs_lo_7 = _bypass_idxs_T_6[1]; // @[CircuitMath.scala 30:8]
  wire [1:0] bypass_idxs_1 = {bypass_idxs_hi_7,bypass_idxs_lo_7}; // @[Cat.scala 30:58]
  wire  bypass_idxs_hi_8 = tail[0]; // @[Lsu.scala 60:12]
  wire [2:0] bypass_idxs_lo_8 = tail[3:1]; // @[Lsu.scala 60:29]
  wire [3:0] _bypass_idxs_T_8 = {bypass_idxs_hi_8,bypass_idxs_lo_8}; // @[Cat.scala 30:58]
  wire [1:0] bypass_idxs_hi_9 = _bypass_idxs_T_8[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] bypass_idxs_lo_9 = _bypass_idxs_T_8[1:0]; // @[OneHot.scala 31:18]
  wire  bypass_idxs_hi_10 = |bypass_idxs_hi_9; // @[OneHot.scala 32:14]
  wire [1:0] _bypass_idxs_T_9 = bypass_idxs_hi_9 | bypass_idxs_lo_9; // @[OneHot.scala 32:28]
  wire  bypass_idxs_lo_10 = _bypass_idxs_T_9[1]; // @[CircuitMath.scala 30:8]
  wire [1:0] bypass_idxs_0 = {bypass_idxs_hi_10,bypass_idxs_lo_10}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_221 = 2'h1 == bypass_idxs_0 ? write_buffer_1_addr : write_buffer_0_addr; // @[Lsu.scala 181:67 Lsu.scala 181:67]
  wire [31:0] _GEN_222 = 2'h2 == bypass_idxs_0 ? write_buffer_2_addr : _GEN_221; // @[Lsu.scala 181:67 Lsu.scala 181:67]
  wire [31:0] _GEN_223 = 2'h3 == bypass_idxs_0 ? write_buffer_3_addr : _GEN_222; // @[Lsu.scala 181:67 Lsu.scala 181:67]
  wire  _GEN_225 = 2'h1 == bypass_idxs_0 ? write_buffer_uncache_1 : write_buffer_uncache_0; // @[Lsu.scala 181:137 Lsu.scala 181:137]
  wire  _GEN_226 = 2'h2 == bypass_idxs_0 ? write_buffer_uncache_2 : _GEN_225; // @[Lsu.scala 181:137 Lsu.scala 181:137]
  wire  _GEN_227 = 2'h3 == bypass_idxs_0 ? write_buffer_uncache_3 : _GEN_226; // @[Lsu.scala 181:137 Lsu.scala 181:137]
  wire  _GEN_229 = 2'h1 == bypass_idxs_0 ? write_buffer_complete_1 : write_buffer_complete_0; // @[Lsu.scala 181:134 Lsu.scala 181:134]
  wire  _GEN_230 = 2'h2 == bypass_idxs_0 ? write_buffer_complete_2 : _GEN_229; // @[Lsu.scala 181:134 Lsu.scala 181:134]
  wire  _GEN_231 = 2'h3 == bypass_idxs_0 ? write_buffer_complete_3 : _GEN_230; // @[Lsu.scala 181:134 Lsu.scala 181:134]
  wire  _GEN_233 = 2'h1 == bypass_idxs_0 ? write_buffer_valid_1 : write_buffer_valid_0; // @[Lsu.scala 181:106 Lsu.scala 181:106]
  wire  _GEN_234 = 2'h2 == bypass_idxs_0 ? write_buffer_valid_2 : _GEN_233; // @[Lsu.scala 181:106 Lsu.scala 181:106]
  wire  _GEN_235 = 2'h3 == bypass_idxs_0 ? write_buffer_valid_3 : _GEN_234; // @[Lsu.scala 181:106 Lsu.scala 181:106]
  wire  hit_buffer_mask_0 = _GEN_223 == mem_addr & (_GEN_235 | _GEN_231 & ~_GEN_227); // @[Lsu.scala 181:80]
  wire [31:0] _GEN_237 = 2'h1 == bypass_idxs_1 ? write_buffer_1_addr : write_buffer_0_addr; // @[Lsu.scala 181:67 Lsu.scala 181:67]
  wire [31:0] _GEN_238 = 2'h2 == bypass_idxs_1 ? write_buffer_2_addr : _GEN_237; // @[Lsu.scala 181:67 Lsu.scala 181:67]
  wire [31:0] _GEN_239 = 2'h3 == bypass_idxs_1 ? write_buffer_3_addr : _GEN_238; // @[Lsu.scala 181:67 Lsu.scala 181:67]
  wire  _GEN_241 = 2'h1 == bypass_idxs_1 ? write_buffer_uncache_1 : write_buffer_uncache_0; // @[Lsu.scala 181:137 Lsu.scala 181:137]
  wire  _GEN_242 = 2'h2 == bypass_idxs_1 ? write_buffer_uncache_2 : _GEN_241; // @[Lsu.scala 181:137 Lsu.scala 181:137]
  wire  _GEN_243 = 2'h3 == bypass_idxs_1 ? write_buffer_uncache_3 : _GEN_242; // @[Lsu.scala 181:137 Lsu.scala 181:137]
  wire  _GEN_245 = 2'h1 == bypass_idxs_1 ? write_buffer_complete_1 : write_buffer_complete_0; // @[Lsu.scala 181:134 Lsu.scala 181:134]
  wire  _GEN_246 = 2'h2 == bypass_idxs_1 ? write_buffer_complete_2 : _GEN_245; // @[Lsu.scala 181:134 Lsu.scala 181:134]
  wire  _GEN_247 = 2'h3 == bypass_idxs_1 ? write_buffer_complete_3 : _GEN_246; // @[Lsu.scala 181:134 Lsu.scala 181:134]
  wire  _GEN_249 = 2'h1 == bypass_idxs_1 ? write_buffer_valid_1 : write_buffer_valid_0; // @[Lsu.scala 181:106 Lsu.scala 181:106]
  wire  _GEN_250 = 2'h2 == bypass_idxs_1 ? write_buffer_valid_2 : _GEN_249; // @[Lsu.scala 181:106 Lsu.scala 181:106]
  wire  _GEN_251 = 2'h3 == bypass_idxs_1 ? write_buffer_valid_3 : _GEN_250; // @[Lsu.scala 181:106 Lsu.scala 181:106]
  wire  hit_buffer_mask_1 = _GEN_239 == mem_addr & (_GEN_251 | _GEN_247 & ~_GEN_243); // @[Lsu.scala 181:80]
  wire [31:0] _GEN_253 = 2'h1 == bypass_idxs_2 ? write_buffer_1_addr : write_buffer_0_addr; // @[Lsu.scala 181:67 Lsu.scala 181:67]
  wire [31:0] _GEN_254 = 2'h2 == bypass_idxs_2 ? write_buffer_2_addr : _GEN_253; // @[Lsu.scala 181:67 Lsu.scala 181:67]
  wire [31:0] _GEN_255 = 2'h3 == bypass_idxs_2 ? write_buffer_3_addr : _GEN_254; // @[Lsu.scala 181:67 Lsu.scala 181:67]
  wire  _GEN_257 = 2'h1 == bypass_idxs_2 ? write_buffer_uncache_1 : write_buffer_uncache_0; // @[Lsu.scala 181:137 Lsu.scala 181:137]
  wire  _GEN_258 = 2'h2 == bypass_idxs_2 ? write_buffer_uncache_2 : _GEN_257; // @[Lsu.scala 181:137 Lsu.scala 181:137]
  wire  _GEN_259 = 2'h3 == bypass_idxs_2 ? write_buffer_uncache_3 : _GEN_258; // @[Lsu.scala 181:137 Lsu.scala 181:137]
  wire  _GEN_261 = 2'h1 == bypass_idxs_2 ? write_buffer_complete_1 : write_buffer_complete_0; // @[Lsu.scala 181:134 Lsu.scala 181:134]
  wire  _GEN_262 = 2'h2 == bypass_idxs_2 ? write_buffer_complete_2 : _GEN_261; // @[Lsu.scala 181:134 Lsu.scala 181:134]
  wire  _GEN_263 = 2'h3 == bypass_idxs_2 ? write_buffer_complete_3 : _GEN_262; // @[Lsu.scala 181:134 Lsu.scala 181:134]
  wire  _GEN_265 = 2'h1 == bypass_idxs_2 ? write_buffer_valid_1 : write_buffer_valid_0; // @[Lsu.scala 181:106 Lsu.scala 181:106]
  wire  _GEN_266 = 2'h2 == bypass_idxs_2 ? write_buffer_valid_2 : _GEN_265; // @[Lsu.scala 181:106 Lsu.scala 181:106]
  wire  _GEN_267 = 2'h3 == bypass_idxs_2 ? write_buffer_valid_3 : _GEN_266; // @[Lsu.scala 181:106 Lsu.scala 181:106]
  wire  hit_buffer_mask_2 = _GEN_255 == mem_addr & (_GEN_267 | _GEN_263 & ~_GEN_259); // @[Lsu.scala 181:80]
  wire [31:0] _GEN_269 = 2'h1 == enq_idx ? write_buffer_1_addr : write_buffer_0_addr; // @[Lsu.scala 181:67 Lsu.scala 181:67]
  wire [31:0] _GEN_270 = 2'h2 == enq_idx ? write_buffer_2_addr : _GEN_269; // @[Lsu.scala 181:67 Lsu.scala 181:67]
  wire [31:0] _GEN_271 = 2'h3 == enq_idx ? write_buffer_3_addr : _GEN_270; // @[Lsu.scala 181:67 Lsu.scala 181:67]
  wire  _GEN_273 = 2'h1 == enq_idx ? write_buffer_uncache_1 : write_buffer_uncache_0; // @[Lsu.scala 181:137 Lsu.scala 181:137]
  wire  _GEN_274 = 2'h2 == enq_idx ? write_buffer_uncache_2 : _GEN_273; // @[Lsu.scala 181:137 Lsu.scala 181:137]
  wire  _GEN_275 = 2'h3 == enq_idx ? write_buffer_uncache_3 : _GEN_274; // @[Lsu.scala 181:137 Lsu.scala 181:137]
  wire  _GEN_277 = 2'h1 == enq_idx ? write_buffer_complete_1 : write_buffer_complete_0; // @[Lsu.scala 181:134 Lsu.scala 181:134]
  wire  _GEN_278 = 2'h2 == enq_idx ? write_buffer_complete_2 : _GEN_277; // @[Lsu.scala 181:134 Lsu.scala 181:134]
  wire  _GEN_279 = 2'h3 == enq_idx ? write_buffer_complete_3 : _GEN_278; // @[Lsu.scala 181:134 Lsu.scala 181:134]
  wire  _GEN_281 = 2'h1 == enq_idx ? write_buffer_valid_1 : write_buffer_valid_0; // @[Lsu.scala 181:106 Lsu.scala 181:106]
  wire  _GEN_282 = 2'h2 == enq_idx ? write_buffer_valid_2 : _GEN_281; // @[Lsu.scala 181:106 Lsu.scala 181:106]
  wire  _GEN_283 = 2'h3 == enq_idx ? write_buffer_valid_3 : _GEN_282; // @[Lsu.scala 181:106 Lsu.scala 181:106]
  wire  hit_buffer_mask_3 = _GEN_271 == mem_addr & (_GEN_283 | _GEN_279 & ~_GEN_275); // @[Lsu.scala 181:80]
  wire [1:0] _hit_buffer_idx_T = hit_buffer_mask_2 ? 2'h2 : 2'h3; // @[Mux.scala 47:69]
  wire [1:0] _hit_buffer_idx_T_1 = hit_buffer_mask_1 ? 2'h1 : _hit_buffer_idx_T; // @[Mux.scala 47:69]
  wire [1:0] _hit_buffer_idx_T_2 = hit_buffer_mask_0 ? 2'h0 : _hit_buffer_idx_T_1; // @[Mux.scala 47:69]
  wire  hit_buffer = hit_buffer_mask_0 | hit_buffer_mask_1 | hit_buffer_mask_2 | hit_buffer_mask_3; // @[Lsu.scala 183:50]
  wire  op_complete = do_enq | do_read & (hit_buffer | io_cache_read_ready); // @[Lsu.scala 186:31]
  wire [1:0] _GEN_285 = 2'h1 == _hit_buffer_idx_T_2 ? bypass_idxs_1 : bypass_idxs_0; // @[Lsu.scala 187:27 Lsu.scala 187:27]
  wire [1:0] _GEN_286 = 2'h2 == _hit_buffer_idx_T_2 ? bypass_idxs_2 : _GEN_285; // @[Lsu.scala 187:27 Lsu.scala 187:27]
  wire [1:0] _GEN_287 = 2'h3 == _hit_buffer_idx_T_2 ? enq_idx : _GEN_286; // @[Lsu.scala 187:27 Lsu.scala 187:27]
  wire [31:0] _GEN_289 = 2'h1 == _GEN_287 ? write_buffer_1_data : write_buffer_0_data; // @[Lsu.scala 187:27 Lsu.scala 187:27]
  wire [31:0] _GEN_290 = 2'h2 == _GEN_287 ? write_buffer_2_data : _GEN_289; // @[Lsu.scala 187:27 Lsu.scala 187:27]
  wire [31:0] _GEN_291 = 2'h3 == _GEN_287 ? write_buffer_3_data : _GEN_290; // @[Lsu.scala 187:27 Lsu.scala 187:27]
  wire [31:0] load_data = hit_buffer ? _GEN_291 : io_cache_resp_data; // @[Lsu.scala 187:27]
  wire  _load_byte_data_T_1 = mem_addr[1:0] == 2'h0; // @[Lsu.scala 188:68]
  wire [7:0] _load_byte_data_T_3 = _load_byte_data_T_1 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _load_byte_data_T_5 = _load_byte_data_T_3 & load_data[7:0]; // @[Lsu.scala 188:82]
  wire  _load_byte_data_T_7 = mem_addr[1:0] == 2'h1; // @[Lsu.scala 188:68]
  wire [7:0] _load_byte_data_T_9 = _load_byte_data_T_7 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _load_byte_data_T_11 = _load_byte_data_T_9 & load_data[15:8]; // @[Lsu.scala 188:82]
  wire  _load_byte_data_T_13 = mem_addr[1:0] == 2'h2; // @[Lsu.scala 188:68]
  wire [7:0] _load_byte_data_T_15 = _load_byte_data_T_13 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _load_byte_data_T_17 = _load_byte_data_T_15 & load_data[23:16]; // @[Lsu.scala 188:82]
  wire  _load_byte_data_T_19 = mem_addr[1:0] == 2'h3; // @[Lsu.scala 188:68]
  wire [7:0] _load_byte_data_T_21 = _load_byte_data_T_19 ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _load_byte_data_T_23 = _load_byte_data_T_21 & load_data[31:24]; // @[Lsu.scala 188:82]
  wire [7:0] _load_byte_data_T_24 = _load_byte_data_T_5 | _load_byte_data_T_11; // @[Lsu.scala 188:122]
  wire [7:0] _load_byte_data_T_25 = _load_byte_data_T_24 | _load_byte_data_T_17; // @[Lsu.scala 188:122]
  wire [7:0] load_byte_data = _load_byte_data_T_25 | _load_byte_data_T_23; // @[Lsu.scala 188:122]
  wire  _load_half_data_T_1 = ~mem_addr[1]; // @[Lsu.scala 189:66]
  wire [15:0] _load_half_data_T_3 = _load_half_data_T_1 ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _load_half_data_T_5 = _load_half_data_T_3 & load_data[15:0]; // @[Lsu.scala 189:80]
  wire [15:0] _load_half_data_T_9 = mem_addr[1] ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12]
  wire [15:0] _load_half_data_T_11 = _load_half_data_T_9 & load_data[31:16]; // @[Lsu.scala 189:80]
  wire [15:0] load_half_data = _load_half_data_T_5 | _load_half_data_T_11; // @[Lsu.scala 189:123]
  wire [23:0] load_final_data_hi = load_byte_data[7] ? 24'hffffff : 24'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _load_final_data_T_4 = {load_final_data_hi,load_byte_data}; // @[Cat.scala 30:58]
  wire [31:0] _load_final_data_T_6 = {24'h0,load_byte_data}; // @[Cat.scala 30:58]
  wire [15:0] load_final_data_hi_2 = load_half_data[15] ? 16'hffff : 16'h0; // @[Bitwise.scala 72:12]
  wire [31:0] _load_final_data_T_10 = {load_final_data_hi_2,load_half_data}; // @[Cat.scala 30:58]
  wire [31:0] _load_final_data_T_12 = {16'h0,load_half_data}; // @[Cat.scala 30:58]
  wire [31:0] _load_final_data_T_14 = 6'h2a == dispatch_info_uop ? _load_final_data_T_4 : load_data; // @[Mux.scala 80:57]
  wire [31:0] _load_final_data_T_16 = 6'h2b == dispatch_info_uop ? _load_final_data_T_6 : _load_final_data_T_14; // @[Mux.scala 80:57]
  wire [31:0] _load_final_data_T_18 = 6'h28 == dispatch_info_uop ? _load_final_data_T_10 : _load_final_data_T_16; // @[Mux.scala 80:57]
  wire  _io_dispatch_info_ready_T_1 = ~dispatch_valid | op_complete; // @[Lsu.scala 212:45]
  assign io_dispatch_info_ready = ~dispatch_valid | op_complete; // @[Lsu.scala 212:45]
  assign io_wb_info_valid = op_complete & dispatch_valid; // @[Lsu.scala 231:34]
  assign io_wb_info_bits_rob_idx = dispatch_info_rob_idx; // @[Lsu.scala 227:26]
  assign io_wb_info_bits_data = 6'h29 == dispatch_info_uop ? _load_final_data_T_12 : _load_final_data_T_18; // @[Mux.scala 80:57]
  assign io_cache_read_valid = ~hit_buffer & do_read; // @[Lsu.scala 207:37]
  assign io_cache_read_bits_addr = $signed(dispatch_info_imm_data) + $signed(dispatch_info_op1_data); // @[Lsu.scala 82:105]
  assign io_cache_read_bits_rob_idx = {{1'd0}, dispatch_info_rob_idx}; // @[Lsu.scala 209:30]
  assign io_cache_write_valid = _GEN_192 & _GEN_196; // @[Lsu.scala 163:47]
  assign io_cache_write_bits_addr = 2'h3 == complete_head_idx ? write_buffer_3_addr : _GEN_203; // @[Lsu.scala 165:28 Lsu.scala 165:28]
  assign io_cache_write_bits_data = 2'h3 == complete_head_idx ? write_buffer_3_data : _GEN_199; // @[Lsu.scala 164:28 Lsu.scala 164:28]
  assign io_cache_write_bits_byte_mask = 2'h3 == complete_head_idx ? write_buffer_3_byte_mask : _GEN_207; // @[Lsu.scala 166:33 Lsu.scala 166:33]
  always @(posedge clock) begin
    if (reset) begin // @[Lsu.scala 255:23]
      dispatch_info_uop <= 6'h0; // @[Rob.scala 142:19]
    end else if (io_need_flush) begin // @[Lsu.scala 238:23]
      dispatch_info_uop <= 6'h0; // @[Rob.scala 142:19]
    end else if (_io_dispatch_info_ready_T_1) begin // @[Lsu.scala 234:40]
      dispatch_info_uop <= io_dispatch_info_bits_uop; // @[Lsu.scala 235:19]
    end
    if (reset) begin // @[Lsu.scala 255:23]
      dispatch_info_rob_idx <= 3'h0; // @[Rob.scala 144:19]
    end else if (io_need_flush) begin // @[Lsu.scala 238:23]
      dispatch_info_rob_idx <= 3'h0; // @[Rob.scala 144:19]
    end else if (_io_dispatch_info_ready_T_1) begin // @[Lsu.scala 234:40]
      dispatch_info_rob_idx <= io_dispatch_info_bits_rob_idx; // @[Lsu.scala 235:19]
    end
    if (reset) begin // @[Lsu.scala 255:23]
      dispatch_info_op1_data <= 32'h0; // @[Rob.scala 146:19]
    end else if (io_need_flush) begin // @[Lsu.scala 238:23]
      dispatch_info_op1_data <= 32'h0; // @[Rob.scala 146:19]
    end else if (_io_dispatch_info_ready_T_1) begin // @[Lsu.scala 234:40]
      dispatch_info_op1_data <= io_dispatch_info_bits_op1_data; // @[Lsu.scala 235:19]
    end
    if (reset) begin // @[Lsu.scala 255:23]
      dispatch_info_op2_data <= 32'h0; // @[Rob.scala 147:19]
    end else if (io_need_flush) begin // @[Lsu.scala 238:23]
      dispatch_info_op2_data <= 32'h0; // @[Rob.scala 147:19]
    end else if (_io_dispatch_info_ready_T_1) begin // @[Lsu.scala 234:40]
      dispatch_info_op2_data <= io_dispatch_info_bits_op2_data; // @[Lsu.scala 235:19]
    end
    if (reset) begin // @[Lsu.scala 255:23]
      dispatch_info_imm_data <= 32'h0; // @[Rob.scala 148:19]
    end else if (io_need_flush) begin // @[Lsu.scala 238:23]
      dispatch_info_imm_data <= 32'h0; // @[Rob.scala 148:19]
    end else if (_io_dispatch_info_ready_T_1) begin // @[Lsu.scala 234:40]
      dispatch_info_imm_data <= io_dispatch_info_bits_imm_data; // @[Lsu.scala 235:19]
    end
    if (reset) begin // @[Lsu.scala 69:38]
      dispatch_valid <= 1'h0; // @[Lsu.scala 69:38]
    end else if (io_need_flush) begin // @[Lsu.scala 238:23]
      dispatch_valid <= 1'h0; // @[Lsu.scala 247:20]
    end else if (_io_dispatch_info_ready_T_1) begin // @[Lsu.scala 234:40]
      dispatch_valid <= io_dispatch_info_valid; // @[Lsu.scala 236:20]
    end
    if (reset) begin // @[Lsu.scala 255:23]
      write_buffer_0_rob_idx <= 4'h0; // @[Lsu.scala 38:15]
    end else if (do_enq) begin // @[Lsu.scala 120:16]
      if (2'h0 == enq_idx) begin // @[Lsu.scala 121:35]
        write_buffer_0_rob_idx <= _write_buffer_enq_idx_rob_idx; // @[Lsu.scala 121:35]
      end
    end
    if (reset) begin // @[Lsu.scala 255:23]
      write_buffer_0_addr <= 32'h0; // @[Lsu.scala 39:15]
    end else if (do_enq) begin // @[Lsu.scala 120:16]
      if (2'h0 == enq_idx) begin // @[Lsu.scala 123:32]
        write_buffer_0_addr <= mem_addr; // @[Lsu.scala 123:32]
      end
    end
    if (reset) begin // @[Lsu.scala 255:23]
      write_buffer_0_data <= 32'h0; // @[Lsu.scala 40:15]
    end else if (do_enq) begin // @[Lsu.scala 120:16]
      if (2'h0 == enq_idx) begin // @[Lsu.scala 122:32]
        write_buffer_0_data <= dispatch_info_op2_data; // @[Lsu.scala 122:32]
      end
    end
    if (reset) begin // @[Lsu.scala 255:23]
      write_buffer_0_byte_mask <= 4'h0; // @[Lsu.scala 41:15]
    end else if (do_enq) begin // @[Lsu.scala 120:16]
      if (2'h0 == enq_idx) begin // @[Lsu.scala 124:37]
        if (6'h24 == dispatch_info_uop) begin // @[Mux.scala 80:57]
          write_buffer_0_byte_mask <= 4'hf;
        end else begin
          write_buffer_0_byte_mask <= _byte_mask_T_22;
        end
      end
    end
    if (reset) begin // @[Lsu.scala 255:23]
      write_buffer_1_rob_idx <= 4'h0; // @[Lsu.scala 38:15]
    end else if (do_enq) begin // @[Lsu.scala 120:16]
      if (2'h1 == enq_idx) begin // @[Lsu.scala 121:35]
        write_buffer_1_rob_idx <= _write_buffer_enq_idx_rob_idx; // @[Lsu.scala 121:35]
      end
    end
    if (reset) begin // @[Lsu.scala 255:23]
      write_buffer_1_addr <= 32'h0; // @[Lsu.scala 39:15]
    end else if (do_enq) begin // @[Lsu.scala 120:16]
      if (2'h1 == enq_idx) begin // @[Lsu.scala 123:32]
        write_buffer_1_addr <= mem_addr; // @[Lsu.scala 123:32]
      end
    end
    if (reset) begin // @[Lsu.scala 255:23]
      write_buffer_1_data <= 32'h0; // @[Lsu.scala 40:15]
    end else if (do_enq) begin // @[Lsu.scala 120:16]
      if (2'h1 == enq_idx) begin // @[Lsu.scala 122:32]
        write_buffer_1_data <= dispatch_info_op2_data; // @[Lsu.scala 122:32]
      end
    end
    if (reset) begin // @[Lsu.scala 255:23]
      write_buffer_1_byte_mask <= 4'h0; // @[Lsu.scala 41:15]
    end else if (do_enq) begin // @[Lsu.scala 120:16]
      if (2'h1 == enq_idx) begin // @[Lsu.scala 124:37]
        if (6'h24 == dispatch_info_uop) begin // @[Mux.scala 80:57]
          write_buffer_1_byte_mask <= 4'hf;
        end else begin
          write_buffer_1_byte_mask <= _byte_mask_T_22;
        end
      end
    end
    if (reset) begin // @[Lsu.scala 255:23]
      write_buffer_2_rob_idx <= 4'h0; // @[Lsu.scala 38:15]
    end else if (do_enq) begin // @[Lsu.scala 120:16]
      if (2'h2 == enq_idx) begin // @[Lsu.scala 121:35]
        write_buffer_2_rob_idx <= _write_buffer_enq_idx_rob_idx; // @[Lsu.scala 121:35]
      end
    end
    if (reset) begin // @[Lsu.scala 255:23]
      write_buffer_2_addr <= 32'h0; // @[Lsu.scala 39:15]
    end else if (do_enq) begin // @[Lsu.scala 120:16]
      if (2'h2 == enq_idx) begin // @[Lsu.scala 123:32]
        write_buffer_2_addr <= mem_addr; // @[Lsu.scala 123:32]
      end
    end
    if (reset) begin // @[Lsu.scala 255:23]
      write_buffer_2_data <= 32'h0; // @[Lsu.scala 40:15]
    end else if (do_enq) begin // @[Lsu.scala 120:16]
      if (2'h2 == enq_idx) begin // @[Lsu.scala 122:32]
        write_buffer_2_data <= dispatch_info_op2_data; // @[Lsu.scala 122:32]
      end
    end
    if (reset) begin // @[Lsu.scala 255:23]
      write_buffer_2_byte_mask <= 4'h0; // @[Lsu.scala 41:15]
    end else if (do_enq) begin // @[Lsu.scala 120:16]
      if (2'h2 == enq_idx) begin // @[Lsu.scala 124:37]
        if (6'h24 == dispatch_info_uop) begin // @[Mux.scala 80:57]
          write_buffer_2_byte_mask <= 4'hf;
        end else begin
          write_buffer_2_byte_mask <= _byte_mask_T_22;
        end
      end
    end
    if (reset) begin // @[Lsu.scala 255:23]
      write_buffer_3_rob_idx <= 4'h0; // @[Lsu.scala 38:15]
    end else if (do_enq) begin // @[Lsu.scala 120:16]
      if (2'h3 == enq_idx) begin // @[Lsu.scala 121:35]
        write_buffer_3_rob_idx <= _write_buffer_enq_idx_rob_idx; // @[Lsu.scala 121:35]
      end
    end
    if (reset) begin // @[Lsu.scala 255:23]
      write_buffer_3_addr <= 32'h0; // @[Lsu.scala 39:15]
    end else if (do_enq) begin // @[Lsu.scala 120:16]
      if (2'h3 == enq_idx) begin // @[Lsu.scala 123:32]
        write_buffer_3_addr <= mem_addr; // @[Lsu.scala 123:32]
      end
    end
    if (reset) begin // @[Lsu.scala 255:23]
      write_buffer_3_data <= 32'h0; // @[Lsu.scala 40:15]
    end else if (do_enq) begin // @[Lsu.scala 120:16]
      if (2'h3 == enq_idx) begin // @[Lsu.scala 122:32]
        write_buffer_3_data <= dispatch_info_op2_data; // @[Lsu.scala 122:32]
      end
    end
    if (reset) begin // @[Lsu.scala 255:23]
      write_buffer_3_byte_mask <= 4'h0; // @[Lsu.scala 41:15]
    end else if (do_enq) begin // @[Lsu.scala 120:16]
      if (2'h3 == enq_idx) begin // @[Lsu.scala 124:37]
        if (6'h24 == dispatch_info_uop) begin // @[Mux.scala 80:57]
          write_buffer_3_byte_mask <= 4'hf;
        end else begin
          write_buffer_3_byte_mask <= _byte_mask_T_22;
        end
      end
    end
    if (reset) begin // @[Lsu.scala 71:38]
      write_buffer_valid_0 <= 1'h0; // @[Lsu.scala 71:38]
    end else if (io_need_flush) begin // @[Lsu.scala 238:23]
      if (~write_buffer_complete_0 & ~will_complete_0) begin // @[Lsu.scala 240:60]
        write_buffer_valid_0 <= 1'h0; // @[Lsu.scala 241:31]
      end else begin
        write_buffer_valid_0 <= _GEN_214;
      end
    end else begin
      write_buffer_valid_0 <= _GEN_214;
    end
    if (reset) begin // @[Lsu.scala 71:38]
      write_buffer_valid_1 <= 1'h0; // @[Lsu.scala 71:38]
    end else if (io_need_flush) begin // @[Lsu.scala 238:23]
      if (~write_buffer_complete_1 & ~will_complete_1) begin // @[Lsu.scala 240:60]
        write_buffer_valid_1 <= 1'h0; // @[Lsu.scala 241:31]
      end else begin
        write_buffer_valid_1 <= _GEN_215;
      end
    end else begin
      write_buffer_valid_1 <= _GEN_215;
    end
    if (reset) begin // @[Lsu.scala 71:38]
      write_buffer_valid_2 <= 1'h0; // @[Lsu.scala 71:38]
    end else if (io_need_flush) begin // @[Lsu.scala 238:23]
      if (~write_buffer_complete_2 & ~will_complete_2) begin // @[Lsu.scala 240:60]
        write_buffer_valid_2 <= 1'h0; // @[Lsu.scala 241:31]
      end else begin
        write_buffer_valid_2 <= _GEN_216;
      end
    end else begin
      write_buffer_valid_2 <= _GEN_216;
    end
    if (reset) begin // @[Lsu.scala 71:38]
      write_buffer_valid_3 <= 1'h0; // @[Lsu.scala 71:38]
    end else if (io_need_flush) begin // @[Lsu.scala 238:23]
      if (~write_buffer_complete_3 & ~will_complete_3) begin // @[Lsu.scala 240:60]
        write_buffer_valid_3 <= 1'h0; // @[Lsu.scala 241:31]
      end else begin
        write_buffer_valid_3 <= _GEN_217;
      end
    end else begin
      write_buffer_valid_3 <= _GEN_217;
    end
    if (reset) begin // @[Lsu.scala 72:38]
      write_buffer_waiting_0 <= 1'h0; // @[Lsu.scala 72:38]
    end else if (io_need_flush) begin // @[Lsu.scala 238:23]
      if (~write_buffer_complete_0 & ~will_complete_0) begin // @[Lsu.scala 240:60]
        write_buffer_waiting_0 <= 1'h0; // @[Lsu.scala 242:33]
      end else begin
        write_buffer_waiting_0 <= _GEN_180;
      end
    end else begin
      write_buffer_waiting_0 <= _GEN_180;
    end
    if (reset) begin // @[Lsu.scala 72:38]
      write_buffer_waiting_1 <= 1'h0; // @[Lsu.scala 72:38]
    end else if (io_need_flush) begin // @[Lsu.scala 238:23]
      if (~write_buffer_complete_1 & ~will_complete_1) begin // @[Lsu.scala 240:60]
        write_buffer_waiting_1 <= 1'h0; // @[Lsu.scala 242:33]
      end else begin
        write_buffer_waiting_1 <= _GEN_181;
      end
    end else begin
      write_buffer_waiting_1 <= _GEN_181;
    end
    if (reset) begin // @[Lsu.scala 72:38]
      write_buffer_waiting_2 <= 1'h0; // @[Lsu.scala 72:38]
    end else if (io_need_flush) begin // @[Lsu.scala 238:23]
      if (~write_buffer_complete_2 & ~will_complete_2) begin // @[Lsu.scala 240:60]
        write_buffer_waiting_2 <= 1'h0; // @[Lsu.scala 242:33]
      end else begin
        write_buffer_waiting_2 <= _GEN_182;
      end
    end else begin
      write_buffer_waiting_2 <= _GEN_182;
    end
    if (reset) begin // @[Lsu.scala 72:38]
      write_buffer_waiting_3 <= 1'h0; // @[Lsu.scala 72:38]
    end else if (io_need_flush) begin // @[Lsu.scala 238:23]
      if (~write_buffer_complete_3 & ~will_complete_3) begin // @[Lsu.scala 240:60]
        write_buffer_waiting_3 <= 1'h0; // @[Lsu.scala 242:33]
      end else begin
        write_buffer_waiting_3 <= _GEN_183;
      end
    end else begin
      write_buffer_waiting_3 <= _GEN_183;
    end
    if (reset) begin // @[Lsu.scala 73:38]
      write_buffer_complete_0 <= 1'h0; // @[Lsu.scala 73:38]
    end else if (_GEN_130 & _GEN_134 & io_rob_commit_1_valid & _GEN_381 == _GEN_138) begin // @[Lsu.scala 142:172]
      write_buffer_complete_0 <= _GEN_164;
    end else if (_GEN_130 & _GEN_134 & io_rob_commit_0_valid & _GEN_376 == _GEN_138) begin // @[Lsu.scala 142:172]
      write_buffer_complete_0 <= _GEN_139;
    end else if (_GEN_68 & _GEN_72 & io_rob_commit_1_valid & _GEN_381 == _GEN_76) begin // @[Lsu.scala 142:172]
      write_buffer_complete_0 <= _GEN_102;
    end else begin
      write_buffer_complete_0 <= _GEN_89;
    end
    if (reset) begin // @[Lsu.scala 73:38]
      write_buffer_complete_1 <= 1'h0; // @[Lsu.scala 73:38]
    end else if (_GEN_130 & _GEN_134 & io_rob_commit_1_valid & _GEN_381 == _GEN_138) begin // @[Lsu.scala 142:172]
      write_buffer_complete_1 <= _GEN_165;
    end else if (_GEN_130 & _GEN_134 & io_rob_commit_0_valid & _GEN_376 == _GEN_138) begin // @[Lsu.scala 142:172]
      write_buffer_complete_1 <= _GEN_140;
    end else if (_GEN_68 & _GEN_72 & io_rob_commit_1_valid & _GEN_381 == _GEN_76) begin // @[Lsu.scala 142:172]
      write_buffer_complete_1 <= _GEN_103;
    end else begin
      write_buffer_complete_1 <= _GEN_90;
    end
    if (reset) begin // @[Lsu.scala 73:38]
      write_buffer_complete_2 <= 1'h0; // @[Lsu.scala 73:38]
    end else if (_GEN_130 & _GEN_134 & io_rob_commit_1_valid & _GEN_381 == _GEN_138) begin // @[Lsu.scala 142:172]
      write_buffer_complete_2 <= _GEN_166;
    end else if (_GEN_130 & _GEN_134 & io_rob_commit_0_valid & _GEN_376 == _GEN_138) begin // @[Lsu.scala 142:172]
      write_buffer_complete_2 <= _GEN_141;
    end else if (_GEN_68 & _GEN_72 & io_rob_commit_1_valid & _GEN_381 == _GEN_76) begin // @[Lsu.scala 142:172]
      write_buffer_complete_2 <= _GEN_104;
    end else begin
      write_buffer_complete_2 <= _GEN_91;
    end
    if (reset) begin // @[Lsu.scala 73:38]
      write_buffer_complete_3 <= 1'h0; // @[Lsu.scala 73:38]
    end else if (_GEN_130 & _GEN_134 & io_rob_commit_1_valid & _GEN_381 == _GEN_138) begin // @[Lsu.scala 142:172]
      write_buffer_complete_3 <= _GEN_167;
    end else if (_GEN_130 & _GEN_134 & io_rob_commit_0_valid & _GEN_376 == _GEN_138) begin // @[Lsu.scala 142:172]
      write_buffer_complete_3 <= _GEN_142;
    end else if (_GEN_68 & _GEN_72 & io_rob_commit_1_valid & _GEN_381 == _GEN_76) begin // @[Lsu.scala 142:172]
      write_buffer_complete_3 <= _GEN_105;
    end else begin
      write_buffer_complete_3 <= _GEN_92;
    end
    if (reset) begin // @[Lsu.scala 74:38]
      write_buffer_uncache_0 <= 1'h0; // @[Lsu.scala 74:38]
    end else if (do_enq) begin // @[Lsu.scala 120:16]
      if (2'h0 == enq_idx) begin // @[Lsu.scala 128:35]
        write_buffer_uncache_0 <= is_uncache; // @[Lsu.scala 128:35]
      end
    end
    if (reset) begin // @[Lsu.scala 74:38]
      write_buffer_uncache_1 <= 1'h0; // @[Lsu.scala 74:38]
    end else if (do_enq) begin // @[Lsu.scala 120:16]
      if (2'h1 == enq_idx) begin // @[Lsu.scala 128:35]
        write_buffer_uncache_1 <= is_uncache; // @[Lsu.scala 128:35]
      end
    end
    if (reset) begin // @[Lsu.scala 74:38]
      write_buffer_uncache_2 <= 1'h0; // @[Lsu.scala 74:38]
    end else if (do_enq) begin // @[Lsu.scala 120:16]
      if (2'h2 == enq_idx) begin // @[Lsu.scala 128:35]
        write_buffer_uncache_2 <= is_uncache; // @[Lsu.scala 128:35]
      end
    end
    if (reset) begin // @[Lsu.scala 74:38]
      write_buffer_uncache_3 <= 1'h0; // @[Lsu.scala 74:38]
    end else if (do_enq) begin // @[Lsu.scala 120:16]
      if (2'h3 == enq_idx) begin // @[Lsu.scala 128:35]
        write_buffer_uncache_3 <= is_uncache; // @[Lsu.scala 128:35]
      end
    end
    if (reset) begin // @[Lsu.scala 75:38]
      complete_head <= 4'h1; // @[Lsu.scala 75:38]
    end else if (io_cache_write_ready) begin // @[Lsu.scala 168:16]
      complete_head <= _complete_head_T; // @[Lsu.scala 169:19]
    end
    if (reset) begin // @[Lsu.scala 76:38]
      tail <= 4'h1; // @[Lsu.scala 76:38]
    end else if (io_need_flush) begin // @[Lsu.scala 238:23]
      if (ready_valid_1 & _T_18 != tail) begin // @[Lsu.scala 152:26]
        tail <= ready_deq_idxs_2;
      end else if (ready_valid_0 & ready_deq_idxs_0 != tail) begin // @[Lsu.scala 152:26]
        tail <= ready_deq_idxs_1;
      end else begin
        tail <= ready_deq_idxs_0;
      end
    end else if (do_enq) begin // @[Lsu.scala 120:16]
      tail <= _tail_T; // @[Lsu.scala 129:10]
    end
    if (reset) begin // @[Lsu.scala 77:38]
      maybe_full <= 1'h0; // @[Lsu.scala 77:38]
    end else if (io_need_flush) begin // @[Lsu.scala 238:23]
      maybe_full <= 1'h0; // @[Lsu.scala 248:16]
    end else begin
      maybe_full <= _GEN_219;
    end
    if (reset) begin // @[Lsu.scala 133:31]
      ready_deq_idxs_0 <= 4'h1; // @[Lsu.scala 133:31]
    end else if (ready_valid_1 & _T_18 != tail) begin // @[Lsu.scala 152:26]
      ready_deq_idxs_0 <= ready_deq_idxs_2;
    end else if (ready_valid_0 & ready_deq_idxs_0 != tail) begin // @[Lsu.scala 152:26]
      ready_deq_idxs_0 <= ready_deq_idxs_1;
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  dispatch_info_uop = _RAND_0[5:0];
  _RAND_1 = {1{`RANDOM}};
  dispatch_info_rob_idx = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  dispatch_info_op1_data = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  dispatch_info_op2_data = _RAND_3[31:0];
  _RAND_4 = {1{`RANDOM}};
  dispatch_info_imm_data = _RAND_4[31:0];
  _RAND_5 = {1{`RANDOM}};
  dispatch_valid = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  write_buffer_0_rob_idx = _RAND_6[3:0];
  _RAND_7 = {1{`RANDOM}};
  write_buffer_0_addr = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  write_buffer_0_data = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  write_buffer_0_byte_mask = _RAND_9[3:0];
  _RAND_10 = {1{`RANDOM}};
  write_buffer_1_rob_idx = _RAND_10[3:0];
  _RAND_11 = {1{`RANDOM}};
  write_buffer_1_addr = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  write_buffer_1_data = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  write_buffer_1_byte_mask = _RAND_13[3:0];
  _RAND_14 = {1{`RANDOM}};
  write_buffer_2_rob_idx = _RAND_14[3:0];
  _RAND_15 = {1{`RANDOM}};
  write_buffer_2_addr = _RAND_15[31:0];
  _RAND_16 = {1{`RANDOM}};
  write_buffer_2_data = _RAND_16[31:0];
  _RAND_17 = {1{`RANDOM}};
  write_buffer_2_byte_mask = _RAND_17[3:0];
  _RAND_18 = {1{`RANDOM}};
  write_buffer_3_rob_idx = _RAND_18[3:0];
  _RAND_19 = {1{`RANDOM}};
  write_buffer_3_addr = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  write_buffer_3_data = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  write_buffer_3_byte_mask = _RAND_21[3:0];
  _RAND_22 = {1{`RANDOM}};
  write_buffer_valid_0 = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  write_buffer_valid_1 = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  write_buffer_valid_2 = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  write_buffer_valid_3 = _RAND_25[0:0];
  _RAND_26 = {1{`RANDOM}};
  write_buffer_waiting_0 = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  write_buffer_waiting_1 = _RAND_27[0:0];
  _RAND_28 = {1{`RANDOM}};
  write_buffer_waiting_2 = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  write_buffer_waiting_3 = _RAND_29[0:0];
  _RAND_30 = {1{`RANDOM}};
  write_buffer_complete_0 = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  write_buffer_complete_1 = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  write_buffer_complete_2 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  write_buffer_complete_3 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  write_buffer_uncache_0 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  write_buffer_uncache_1 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  write_buffer_uncache_2 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  write_buffer_uncache_3 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  complete_head = _RAND_38[3:0];
  _RAND_39 = {1{`RANDOM}};
  tail = _RAND_39[3:0];
  _RAND_40 = {1{`RANDOM}};
  maybe_full = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  ready_deq_idxs_0 = _RAND_41[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Mdu(
  input         clock,
  input         reset,
  input         io_dispatch_info_valid,
  input  [2:0]  io_dispatch_info_bits_rob_idx,
  input  [31:0] io_dispatch_info_bits_op1_data,
  input  [31:0] io_dispatch_info_bits_op2_data,
  output        io_wb_info_valid,
  output [2:0]  io_wb_info_bits_rob_idx,
  output [31:0] io_wb_info_bits_data,
  input         io_need_flush
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] dispatch_info_rob_idx; // @[Mdu.scala 20:34]
  reg [31:0] dispatch_info_op1_data; // @[Mdu.scala 20:34]
  reg [31:0] dispatch_info_op2_data; // @[Mdu.scala 20:34]
  reg  dispatch_valid; // @[Mdu.scala 22:38]
  wire [63:0] result = dispatch_info_op1_data * dispatch_info_op2_data; // @[Mdu.scala 26:38]
  assign io_wb_info_valid = dispatch_valid; // @[Mdu.scala 47:19]
  assign io_wb_info_bits_rob_idx = dispatch_info_rob_idx; // @[Mdu.scala 43:26]
  assign io_wb_info_bits_data = result[31:0]; // @[Mdu.scala 42:31]
  always @(posedge clock) begin
    if (reset) begin // @[Mdu.scala 56:23]
      dispatch_info_rob_idx <= 3'h0; // @[Rob.scala 144:19]
    end else if (io_need_flush) begin // @[Mdu.scala 49:22]
      dispatch_info_rob_idx <= 3'h0; // @[Rob.scala 144:19]
    end else begin
      dispatch_info_rob_idx <= io_dispatch_info_bits_rob_idx; // @[Mdu.scala 21:17]
    end
    if (reset) begin // @[Mdu.scala 56:23]
      dispatch_info_op1_data <= 32'h0; // @[Rob.scala 146:19]
    end else if (io_need_flush) begin // @[Mdu.scala 49:22]
      dispatch_info_op1_data <= 32'h0; // @[Rob.scala 146:19]
    end else begin
      dispatch_info_op1_data <= io_dispatch_info_bits_op1_data; // @[Mdu.scala 21:17]
    end
    if (reset) begin // @[Mdu.scala 56:23]
      dispatch_info_op2_data <= 32'h0; // @[Rob.scala 147:19]
    end else if (io_need_flush) begin // @[Mdu.scala 49:22]
      dispatch_info_op2_data <= 32'h0; // @[Rob.scala 147:19]
    end else begin
      dispatch_info_op2_data <= io_dispatch_info_bits_op2_data; // @[Mdu.scala 21:17]
    end
    if (reset) begin // @[Mdu.scala 22:38]
      dispatch_valid <= 1'h0; // @[Mdu.scala 22:38]
    end else if (io_need_flush) begin // @[Mdu.scala 49:22]
      dispatch_valid <= 1'h0; // @[Mdu.scala 51:19]
    end else begin
      dispatch_valid <= io_dispatch_info_valid; // @[Mdu.scala 23:17]
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  dispatch_info_rob_idx = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  dispatch_info_op1_data = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  dispatch_info_op2_data = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  dispatch_valid = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Dcache(
  output        io_dcache_read_req_ready,
  input         io_dcache_read_req_valid,
  input  [31:0] io_dcache_read_req_bits_addr,
  input  [3:0]  io_dcache_read_req_bits_rob_idx,
  output [31:0] io_dcache_read_resp_data,
  output        io_dcache_write_req_ready,
  input         io_dcache_write_req_valid,
  input  [31:0] io_dcache_write_req_bits_addr,
  input  [31:0] io_dcache_write_req_bits_data,
  input  [3:0]  io_dcache_write_req_bits_byte_mask,
  input         io_io_read_req_ready,
  output        io_io_read_req_valid,
  output [31:0] io_io_read_req_bits_addr,
  output [3:0]  io_io_read_req_bits_rob_idx,
  input  [31:0] io_io_read_resp_bits_data,
  input         io_io_write_req_ready,
  output        io_io_write_req_valid,
  output [31:0] io_io_write_req_bits_addr,
  output [31:0] io_io_write_req_bits_data,
  output [3:0]  io_io_write_req_bits_byte_mask
);
  assign io_dcache_read_req_ready = io_io_read_req_ready; // @[Dcache.scala 21:17]
  assign io_dcache_read_resp_data = io_io_read_resp_bits_data; // @[Dcache.scala 22:23]
  assign io_dcache_write_req_ready = io_io_write_req_ready; // @[Dcache.scala 24:18]
  assign io_io_read_req_valid = io_dcache_read_req_valid; // @[Dcache.scala 21:17]
  assign io_io_read_req_bits_addr = io_dcache_read_req_bits_addr; // @[Dcache.scala 21:17]
  assign io_io_read_req_bits_rob_idx = io_dcache_read_req_bits_rob_idx; // @[Dcache.scala 21:17]
  assign io_io_write_req_valid = io_dcache_write_req_valid; // @[Dcache.scala 24:18]
  assign io_io_write_req_bits_addr = io_dcache_write_req_bits_addr; // @[Dcache.scala 24:18]
  assign io_io_write_req_bits_data = io_dcache_write_req_bits_data; // @[Dcache.scala 24:18]
  assign io_io_write_req_bits_byte_mask = io_dcache_write_req_bits_byte_mask; // @[Dcache.scala 24:18]
endmodule
module Exu(
  input         clock,
  input         reset,
  input         io_fb_inst_bank_i_valid,
  input  [31:0] io_fb_inst_bank_i_bits_data_0_inst,
  input  [31:0] io_fb_inst_bank_i_bits_data_0_inst_addr,
  input  [3:0]  io_fb_inst_bank_i_bits_data_0_gh_backup,
  input         io_fb_inst_bank_i_bits_data_0_is_valid,
  input         io_fb_inst_bank_i_bits_data_0_predict_taken,
  input  [31:0] io_fb_inst_bank_i_bits_data_1_inst,
  input  [31:0] io_fb_inst_bank_i_bits_data_1_inst_addr,
  input  [3:0]  io_fb_inst_bank_i_bits_data_1_gh_backup,
  input         io_fb_inst_bank_i_bits_data_1_is_valid,
  input         io_fb_inst_bank_i_bits_data_1_predict_taken,
  output        io_fb_resp_deq_valid_0,
  output        io_fb_resp_deq_valid_1,
  output        io_ex_branch_info_o_valid,
  output [31:0] io_ex_branch_info_o_bits_target_addr,
  output [31:0] io_ex_branch_info_o_bits_inst_addr,
  output [3:0]  io_ex_branch_info_o_bits_gh_update,
  output        io_ex_branch_info_o_bits_is_branch,
  output        io_ex_branch_info_o_bits_is_taken,
  output        io_ex_branch_info_o_bits_predict_miss,
  input         io_dcache_io_read_req_ready,
  output        io_dcache_io_read_req_valid,
  output [31:0] io_dcache_io_read_req_bits_addr,
  output [3:0]  io_dcache_io_read_req_bits_rob_idx,
  input  [31:0] io_dcache_io_read_resp_bits_data,
  input         io_dcache_io_write_req_ready,
  output        io_dcache_io_write_req_valid,
  output [31:0] io_dcache_io_write_req_bits_addr,
  output [31:0] io_dcache_io_write_req_bits_data,
  output [3:0]  io_dcache_io_write_req_bits_byte_mask,
  output        io_need_flush,
  output        io_rob_commit_0_valid,
  output [2:0]  io_rob_commit_0_bits_des_rob,
  output        io_rob_commit_1_valid,
  output [2:0]  io_rob_commit_1_bits_des_rob
);
  wire  decode_clock; // @[Exu.scala 24:22]
  wire  decode_reset; // @[Exu.scala 24:22]
  wire  decode_io_fb_inst_bank_valid; // @[Exu.scala 24:22]
  wire [31:0] decode_io_fb_inst_bank_bits_data_0_inst; // @[Exu.scala 24:22]
  wire [31:0] decode_io_fb_inst_bank_bits_data_0_inst_addr; // @[Exu.scala 24:22]
  wire [3:0] decode_io_fb_inst_bank_bits_data_0_gh_backup; // @[Exu.scala 24:22]
  wire  decode_io_fb_inst_bank_bits_data_0_is_valid; // @[Exu.scala 24:22]
  wire  decode_io_fb_inst_bank_bits_data_0_predict_taken; // @[Exu.scala 24:22]
  wire [31:0] decode_io_fb_inst_bank_bits_data_1_inst; // @[Exu.scala 24:22]
  wire [31:0] decode_io_fb_inst_bank_bits_data_1_inst_addr; // @[Exu.scala 24:22]
  wire [3:0] decode_io_fb_inst_bank_bits_data_1_gh_backup; // @[Exu.scala 24:22]
  wire  decode_io_fb_inst_bank_bits_data_1_is_valid; // @[Exu.scala 24:22]
  wire  decode_io_fb_inst_bank_bits_data_1_predict_taken; // @[Exu.scala 24:22]
  wire  decode_io_fb_resp_deq_valid_0; // @[Exu.scala 24:22]
  wire  decode_io_fb_resp_deq_valid_1; // @[Exu.scala 24:22]
  wire  decode_io_rob_allocate_allocate_req_valid; // @[Exu.scala 24:22]
  wire  decode_io_rob_allocate_allocate_req_bits_0; // @[Exu.scala 24:22]
  wire  decode_io_rob_allocate_allocate_req_bits_1; // @[Exu.scala 24:22]
  wire  decode_io_rob_allocate_allocate_info_valid; // @[Exu.scala 24:22]
  wire [2:0] decode_io_rob_allocate_allocate_info_bits_0_rob_idx; // @[Exu.scala 24:22]
  wire  decode_io_rob_allocate_allocate_info_bits_0_inst_valid; // @[Exu.scala 24:22]
  wire [31:0] decode_io_rob_allocate_allocate_info_bits_0_inst_addr; // @[Exu.scala 24:22]
  wire [5:0] decode_io_rob_allocate_allocate_info_bits_0_uop; // @[Exu.scala 24:22]
  wire [2:0] decode_io_rob_allocate_allocate_info_bits_0_unit_sel; // @[Exu.scala 24:22]
  wire  decode_io_rob_allocate_allocate_info_bits_0_need_imm; // @[Exu.scala 24:22]
  wire [31:0] decode_io_rob_allocate_allocate_info_bits_0_commit_addr; // @[Exu.scala 24:22]
  wire [3:0] decode_io_rob_allocate_allocate_info_bits_0_gh_info; // @[Exu.scala 24:22]
  wire [31:0] decode_io_rob_allocate_allocate_info_bits_0_imm_data; // @[Exu.scala 24:22]
  wire  decode_io_rob_allocate_allocate_info_bits_0_flush_on_commit; // @[Exu.scala 24:22]
  wire  decode_io_rob_allocate_allocate_info_bits_0_predict_taken; // @[Exu.scala 24:22]
  wire [2:0] decode_io_rob_allocate_allocate_info_bits_1_rob_idx; // @[Exu.scala 24:22]
  wire  decode_io_rob_allocate_allocate_info_bits_1_inst_valid; // @[Exu.scala 24:22]
  wire [31:0] decode_io_rob_allocate_allocate_info_bits_1_inst_addr; // @[Exu.scala 24:22]
  wire [5:0] decode_io_rob_allocate_allocate_info_bits_1_uop; // @[Exu.scala 24:22]
  wire [2:0] decode_io_rob_allocate_allocate_info_bits_1_unit_sel; // @[Exu.scala 24:22]
  wire  decode_io_rob_allocate_allocate_info_bits_1_need_imm; // @[Exu.scala 24:22]
  wire [31:0] decode_io_rob_allocate_allocate_info_bits_1_commit_addr; // @[Exu.scala 24:22]
  wire [3:0] decode_io_rob_allocate_allocate_info_bits_1_gh_info; // @[Exu.scala 24:22]
  wire [31:0] decode_io_rob_allocate_allocate_info_bits_1_imm_data; // @[Exu.scala 24:22]
  wire  decode_io_rob_allocate_allocate_info_bits_1_flush_on_commit; // @[Exu.scala 24:22]
  wire  decode_io_rob_allocate_allocate_info_bits_1_predict_taken; // @[Exu.scala 24:22]
  wire  decode_io_rob_allocate_allocate_resp_valid; // @[Exu.scala 24:22]
  wire [2:0] decode_io_rob_allocate_allocate_resp_bits_rob_idx_0; // @[Exu.scala 24:22]
  wire [2:0] decode_io_rob_allocate_allocate_resp_bits_rob_idx_1; // @[Exu.scala 24:22]
  wire  decode_io_rob_allocate_allocate_resp_bits_enq_valid_mask_0; // @[Exu.scala 24:22]
  wire  decode_io_rob_allocate_allocate_resp_bits_enq_valid_mask_1; // @[Exu.scala 24:22]
  wire  decode_io_rename_info_valid; // @[Exu.scala 24:22]
  wire  decode_io_rename_info_bits_0_is_valid; // @[Exu.scala 24:22]
  wire [4:0] decode_io_rename_info_bits_0_op1_addr; // @[Exu.scala 24:22]
  wire [4:0] decode_io_rename_info_bits_0_op2_addr; // @[Exu.scala 24:22]
  wire [4:0] decode_io_rename_info_bits_0_des_addr; // @[Exu.scala 24:22]
  wire [2:0] decode_io_rename_info_bits_0_des_rob; // @[Exu.scala 24:22]
  wire  decode_io_rename_info_bits_1_is_valid; // @[Exu.scala 24:22]
  wire [4:0] decode_io_rename_info_bits_1_op1_addr; // @[Exu.scala 24:22]
  wire [4:0] decode_io_rename_info_bits_1_op2_addr; // @[Exu.scala 24:22]
  wire [4:0] decode_io_rename_info_bits_1_des_addr; // @[Exu.scala 24:22]
  wire [2:0] decode_io_rename_info_bits_1_des_rob; // @[Exu.scala 24:22]
  wire  decode_io_need_flush; // @[Exu.scala 24:22]
  wire  rename_clock; // @[Exu.scala 25:22]
  wire  rename_reset; // @[Exu.scala 25:22]
  wire  rename_io_rename_info_valid; // @[Exu.scala 25:22]
  wire  rename_io_rename_info_bits_0_is_valid; // @[Exu.scala 25:22]
  wire [4:0] rename_io_rename_info_bits_0_op1_addr; // @[Exu.scala 25:22]
  wire [4:0] rename_io_rename_info_bits_0_op2_addr; // @[Exu.scala 25:22]
  wire [4:0] rename_io_rename_info_bits_0_des_addr; // @[Exu.scala 25:22]
  wire [2:0] rename_io_rename_info_bits_0_des_rob; // @[Exu.scala 25:22]
  wire  rename_io_rename_info_bits_1_is_valid; // @[Exu.scala 25:22]
  wire [4:0] rename_io_rename_info_bits_1_op1_addr; // @[Exu.scala 25:22]
  wire [4:0] rename_io_rename_info_bits_1_op2_addr; // @[Exu.scala 25:22]
  wire [4:0] rename_io_rename_info_bits_1_des_addr; // @[Exu.scala 25:22]
  wire [2:0] rename_io_rename_info_bits_1_des_rob; // @[Exu.scala 25:22]
  wire  rename_io_rob_commit_0_valid; // @[Exu.scala 25:22]
  wire [2:0] rename_io_rob_commit_0_bits_des_rob; // @[Exu.scala 25:22]
  wire [4:0] rename_io_rob_commit_0_bits_commit_addr; // @[Exu.scala 25:22]
  wire  rename_io_rob_commit_1_valid; // @[Exu.scala 25:22]
  wire [2:0] rename_io_rob_commit_1_bits_des_rob; // @[Exu.scala 25:22]
  wire [4:0] rename_io_rob_commit_1_bits_commit_addr; // @[Exu.scala 25:22]
  wire [4:0] rename_io_reg_read_0_op1_addr; // @[Exu.scala 25:22]
  wire [4:0] rename_io_reg_read_0_op2_addr; // @[Exu.scala 25:22]
  wire [31:0] rename_io_reg_read_0_op1_data; // @[Exu.scala 25:22]
  wire [31:0] rename_io_reg_read_0_op2_data; // @[Exu.scala 25:22]
  wire [4:0] rename_io_reg_read_1_op1_addr; // @[Exu.scala 25:22]
  wire [4:0] rename_io_reg_read_1_op2_addr; // @[Exu.scala 25:22]
  wire [31:0] rename_io_reg_read_1_op1_data; // @[Exu.scala 25:22]
  wire [31:0] rename_io_reg_read_1_op2_data; // @[Exu.scala 25:22]
  wire  rename_io_rob_init_info_valid; // @[Exu.scala 25:22]
  wire  rename_io_rob_init_info_bits_0_is_valid; // @[Exu.scala 25:22]
  wire [2:0] rename_io_rob_init_info_bits_0_des_rob; // @[Exu.scala 25:22]
  wire [2:0] rename_io_rob_init_info_bits_0_op1_rob; // @[Exu.scala 25:22]
  wire [2:0] rename_io_rob_init_info_bits_0_op2_rob; // @[Exu.scala 25:22]
  wire [31:0] rename_io_rob_init_info_bits_0_op1_regData; // @[Exu.scala 25:22]
  wire [31:0] rename_io_rob_init_info_bits_0_op2_regData; // @[Exu.scala 25:22]
  wire  rename_io_rob_init_info_bits_0_op1_in_rob; // @[Exu.scala 25:22]
  wire  rename_io_rob_init_info_bits_0_op2_in_rob; // @[Exu.scala 25:22]
  wire  rename_io_rob_init_info_bits_1_is_valid; // @[Exu.scala 25:22]
  wire [2:0] rename_io_rob_init_info_bits_1_des_rob; // @[Exu.scala 25:22]
  wire [2:0] rename_io_rob_init_info_bits_1_op1_rob; // @[Exu.scala 25:22]
  wire [2:0] rename_io_rob_init_info_bits_1_op2_rob; // @[Exu.scala 25:22]
  wire [31:0] rename_io_rob_init_info_bits_1_op1_regData; // @[Exu.scala 25:22]
  wire [31:0] rename_io_rob_init_info_bits_1_op2_regData; // @[Exu.scala 25:22]
  wire  rename_io_rob_init_info_bits_1_op1_in_rob; // @[Exu.scala 25:22]
  wire  rename_io_rob_init_info_bits_1_op2_in_rob; // @[Exu.scala 25:22]
  wire  rename_io_need_flush; // @[Exu.scala 25:22]
  wire  regfile_clock; // @[Exu.scala 26:23]
  wire  regfile_reset; // @[Exu.scala 26:23]
  wire [4:0] regfile_io_reg_read_0_op1_addr; // @[Exu.scala 26:23]
  wire [4:0] regfile_io_reg_read_0_op2_addr; // @[Exu.scala 26:23]
  wire [31:0] regfile_io_reg_read_0_op1_data; // @[Exu.scala 26:23]
  wire [31:0] regfile_io_reg_read_0_op2_data; // @[Exu.scala 26:23]
  wire [4:0] regfile_io_reg_read_1_op1_addr; // @[Exu.scala 26:23]
  wire [4:0] regfile_io_reg_read_1_op2_addr; // @[Exu.scala 26:23]
  wire [31:0] regfile_io_reg_read_1_op1_data; // @[Exu.scala 26:23]
  wire [31:0] regfile_io_reg_read_1_op2_data; // @[Exu.scala 26:23]
  wire  regfile_io_rob_commit_i_0_valid; // @[Exu.scala 26:23]
  wire [4:0] regfile_io_rob_commit_i_0_bits_commit_addr; // @[Exu.scala 26:23]
  wire [31:0] regfile_io_rob_commit_i_0_bits_commit_data; // @[Exu.scala 26:23]
  wire  regfile_io_rob_commit_i_1_valid; // @[Exu.scala 26:23]
  wire [4:0] regfile_io_rob_commit_i_1_bits_commit_addr; // @[Exu.scala 26:23]
  wire [31:0] regfile_io_rob_commit_i_1_bits_commit_data; // @[Exu.scala 26:23]
  wire  rob_clock; // @[Exu.scala 27:19]
  wire  rob_reset; // @[Exu.scala 27:19]
  wire  rob_io_rob_allocate_allocate_req_valid; // @[Exu.scala 27:19]
  wire  rob_io_rob_allocate_allocate_req_bits_0; // @[Exu.scala 27:19]
  wire  rob_io_rob_allocate_allocate_req_bits_1; // @[Exu.scala 27:19]
  wire  rob_io_rob_allocate_allocate_info_valid; // @[Exu.scala 27:19]
  wire [2:0] rob_io_rob_allocate_allocate_info_bits_0_rob_idx; // @[Exu.scala 27:19]
  wire  rob_io_rob_allocate_allocate_info_bits_0_inst_valid; // @[Exu.scala 27:19]
  wire [31:0] rob_io_rob_allocate_allocate_info_bits_0_inst_addr; // @[Exu.scala 27:19]
  wire [5:0] rob_io_rob_allocate_allocate_info_bits_0_uop; // @[Exu.scala 27:19]
  wire [2:0] rob_io_rob_allocate_allocate_info_bits_0_unit_sel; // @[Exu.scala 27:19]
  wire  rob_io_rob_allocate_allocate_info_bits_0_need_imm; // @[Exu.scala 27:19]
  wire [31:0] rob_io_rob_allocate_allocate_info_bits_0_commit_addr; // @[Exu.scala 27:19]
  wire [3:0] rob_io_rob_allocate_allocate_info_bits_0_gh_info; // @[Exu.scala 27:19]
  wire [31:0] rob_io_rob_allocate_allocate_info_bits_0_imm_data; // @[Exu.scala 27:19]
  wire  rob_io_rob_allocate_allocate_info_bits_0_flush_on_commit; // @[Exu.scala 27:19]
  wire  rob_io_rob_allocate_allocate_info_bits_0_predict_taken; // @[Exu.scala 27:19]
  wire [2:0] rob_io_rob_allocate_allocate_info_bits_1_rob_idx; // @[Exu.scala 27:19]
  wire  rob_io_rob_allocate_allocate_info_bits_1_inst_valid; // @[Exu.scala 27:19]
  wire [31:0] rob_io_rob_allocate_allocate_info_bits_1_inst_addr; // @[Exu.scala 27:19]
  wire [5:0] rob_io_rob_allocate_allocate_info_bits_1_uop; // @[Exu.scala 27:19]
  wire [2:0] rob_io_rob_allocate_allocate_info_bits_1_unit_sel; // @[Exu.scala 27:19]
  wire  rob_io_rob_allocate_allocate_info_bits_1_need_imm; // @[Exu.scala 27:19]
  wire [31:0] rob_io_rob_allocate_allocate_info_bits_1_commit_addr; // @[Exu.scala 27:19]
  wire [3:0] rob_io_rob_allocate_allocate_info_bits_1_gh_info; // @[Exu.scala 27:19]
  wire [31:0] rob_io_rob_allocate_allocate_info_bits_1_imm_data; // @[Exu.scala 27:19]
  wire  rob_io_rob_allocate_allocate_info_bits_1_flush_on_commit; // @[Exu.scala 27:19]
  wire  rob_io_rob_allocate_allocate_info_bits_1_predict_taken; // @[Exu.scala 27:19]
  wire  rob_io_rob_allocate_allocate_resp_valid; // @[Exu.scala 27:19]
  wire [2:0] rob_io_rob_allocate_allocate_resp_bits_rob_idx_0; // @[Exu.scala 27:19]
  wire [2:0] rob_io_rob_allocate_allocate_resp_bits_rob_idx_1; // @[Exu.scala 27:19]
  wire  rob_io_rob_allocate_allocate_resp_bits_enq_valid_mask_0; // @[Exu.scala 27:19]
  wire  rob_io_rob_allocate_allocate_resp_bits_enq_valid_mask_1; // @[Exu.scala 27:19]
  wire  rob_io_rob_init_info_valid; // @[Exu.scala 27:19]
  wire  rob_io_rob_init_info_bits_0_is_valid; // @[Exu.scala 27:19]
  wire [2:0] rob_io_rob_init_info_bits_0_des_rob; // @[Exu.scala 27:19]
  wire [2:0] rob_io_rob_init_info_bits_0_op1_rob; // @[Exu.scala 27:19]
  wire [2:0] rob_io_rob_init_info_bits_0_op2_rob; // @[Exu.scala 27:19]
  wire [31:0] rob_io_rob_init_info_bits_0_op1_regData; // @[Exu.scala 27:19]
  wire [31:0] rob_io_rob_init_info_bits_0_op2_regData; // @[Exu.scala 27:19]
  wire  rob_io_rob_init_info_bits_0_op1_in_rob; // @[Exu.scala 27:19]
  wire  rob_io_rob_init_info_bits_0_op2_in_rob; // @[Exu.scala 27:19]
  wire  rob_io_rob_init_info_bits_1_is_valid; // @[Exu.scala 27:19]
  wire [2:0] rob_io_rob_init_info_bits_1_des_rob; // @[Exu.scala 27:19]
  wire [2:0] rob_io_rob_init_info_bits_1_op1_rob; // @[Exu.scala 27:19]
  wire [2:0] rob_io_rob_init_info_bits_1_op2_rob; // @[Exu.scala 27:19]
  wire [31:0] rob_io_rob_init_info_bits_1_op1_regData; // @[Exu.scala 27:19]
  wire [31:0] rob_io_rob_init_info_bits_1_op2_regData; // @[Exu.scala 27:19]
  wire  rob_io_rob_init_info_bits_1_op1_in_rob; // @[Exu.scala 27:19]
  wire  rob_io_rob_init_info_bits_1_op2_in_rob; // @[Exu.scala 27:19]
  wire  rob_io_wb_info_i_0_valid; // @[Exu.scala 27:19]
  wire [2:0] rob_io_wb_info_i_0_bits_rob_idx; // @[Exu.scala 27:19]
  wire [31:0] rob_io_wb_info_i_0_bits_data; // @[Exu.scala 27:19]
  wire  rob_io_wb_info_i_1_valid; // @[Exu.scala 27:19]
  wire [2:0] rob_io_wb_info_i_1_bits_rob_idx; // @[Exu.scala 27:19]
  wire [31:0] rob_io_wb_info_i_1_bits_data; // @[Exu.scala 27:19]
  wire  rob_io_wb_info_i_2_valid; // @[Exu.scala 27:19]
  wire [2:0] rob_io_wb_info_i_2_bits_rob_idx; // @[Exu.scala 27:19]
  wire [31:0] rob_io_wb_info_i_2_bits_data; // @[Exu.scala 27:19]
  wire [31:0] rob_io_wb_info_i_2_bits_target_addr; // @[Exu.scala 27:19]
  wire  rob_io_wb_info_i_2_bits_is_taken; // @[Exu.scala 27:19]
  wire  rob_io_wb_info_i_2_bits_predict_miss; // @[Exu.scala 27:19]
  wire  rob_io_wb_info_i_3_valid; // @[Exu.scala 27:19]
  wire [2:0] rob_io_wb_info_i_3_bits_rob_idx; // @[Exu.scala 27:19]
  wire [31:0] rob_io_wb_info_i_3_bits_data; // @[Exu.scala 27:19]
  wire  rob_io_wb_info_i_4_valid; // @[Exu.scala 27:19]
  wire [2:0] rob_io_wb_info_i_4_bits_rob_idx; // @[Exu.scala 27:19]
  wire [31:0] rob_io_wb_info_i_4_bits_data; // @[Exu.scala 27:19]
  wire  rob_io_dispatch_info_o_0_valid; // @[Exu.scala 27:19]
  wire [5:0] rob_io_dispatch_info_o_0_bits_uop; // @[Exu.scala 27:19]
  wire  rob_io_dispatch_info_o_0_bits_need_imm; // @[Exu.scala 27:19]
  wire [2:0] rob_io_dispatch_info_o_0_bits_rob_idx; // @[Exu.scala 27:19]
  wire [31:0] rob_io_dispatch_info_o_0_bits_op1_data; // @[Exu.scala 27:19]
  wire [31:0] rob_io_dispatch_info_o_0_bits_op2_data; // @[Exu.scala 27:19]
  wire [31:0] rob_io_dispatch_info_o_0_bits_imm_data; // @[Exu.scala 27:19]
  wire  rob_io_dispatch_info_o_1_valid; // @[Exu.scala 27:19]
  wire [5:0] rob_io_dispatch_info_o_1_bits_uop; // @[Exu.scala 27:19]
  wire  rob_io_dispatch_info_o_1_bits_need_imm; // @[Exu.scala 27:19]
  wire [2:0] rob_io_dispatch_info_o_1_bits_rob_idx; // @[Exu.scala 27:19]
  wire [31:0] rob_io_dispatch_info_o_1_bits_op1_data; // @[Exu.scala 27:19]
  wire [31:0] rob_io_dispatch_info_o_1_bits_op2_data; // @[Exu.scala 27:19]
  wire [31:0] rob_io_dispatch_info_o_1_bits_imm_data; // @[Exu.scala 27:19]
  wire  rob_io_dispatch_info_o_2_valid; // @[Exu.scala 27:19]
  wire [5:0] rob_io_dispatch_info_o_2_bits_uop; // @[Exu.scala 27:19]
  wire [2:0] rob_io_dispatch_info_o_2_bits_rob_idx; // @[Exu.scala 27:19]
  wire [31:0] rob_io_dispatch_info_o_2_bits_inst_addr; // @[Exu.scala 27:19]
  wire [31:0] rob_io_dispatch_info_o_2_bits_op1_data; // @[Exu.scala 27:19]
  wire [31:0] rob_io_dispatch_info_o_2_bits_op2_data; // @[Exu.scala 27:19]
  wire [31:0] rob_io_dispatch_info_o_2_bits_imm_data; // @[Exu.scala 27:19]
  wire  rob_io_dispatch_info_o_2_bits_predict_taken; // @[Exu.scala 27:19]
  wire  rob_io_dispatch_info_o_3_valid; // @[Exu.scala 27:19]
  wire [2:0] rob_io_dispatch_info_o_3_bits_rob_idx; // @[Exu.scala 27:19]
  wire [31:0] rob_io_dispatch_info_o_3_bits_op1_data; // @[Exu.scala 27:19]
  wire [31:0] rob_io_dispatch_info_o_3_bits_op2_data; // @[Exu.scala 27:19]
  wire  rob_io_dispatch_info_o_4_ready; // @[Exu.scala 27:19]
  wire  rob_io_dispatch_info_o_4_valid; // @[Exu.scala 27:19]
  wire [5:0] rob_io_dispatch_info_o_4_bits_uop; // @[Exu.scala 27:19]
  wire [2:0] rob_io_dispatch_info_o_4_bits_rob_idx; // @[Exu.scala 27:19]
  wire [31:0] rob_io_dispatch_info_o_4_bits_op1_data; // @[Exu.scala 27:19]
  wire [31:0] rob_io_dispatch_info_o_4_bits_op2_data; // @[Exu.scala 27:19]
  wire [31:0] rob_io_dispatch_info_o_4_bits_imm_data; // @[Exu.scala 27:19]
  wire  rob_io_rob_commit_0_valid; // @[Exu.scala 27:19]
  wire [2:0] rob_io_rob_commit_0_bits_des_rob; // @[Exu.scala 27:19]
  wire [4:0] rob_io_rob_commit_0_bits_commit_addr; // @[Exu.scala 27:19]
  wire [31:0] rob_io_rob_commit_0_bits_commit_data; // @[Exu.scala 27:19]
  wire  rob_io_rob_commit_1_valid; // @[Exu.scala 27:19]
  wire [2:0] rob_io_rob_commit_1_bits_des_rob; // @[Exu.scala 27:19]
  wire [4:0] rob_io_rob_commit_1_bits_commit_addr; // @[Exu.scala 27:19]
  wire [31:0] rob_io_rob_commit_1_bits_commit_data; // @[Exu.scala 27:19]
  wire  rob_io_branch_info_valid; // @[Exu.scala 27:19]
  wire [31:0] rob_io_branch_info_bits_target_addr; // @[Exu.scala 27:19]
  wire [31:0] rob_io_branch_info_bits_inst_addr; // @[Exu.scala 27:19]
  wire [3:0] rob_io_branch_info_bits_gh_update; // @[Exu.scala 27:19]
  wire  rob_io_branch_info_bits_is_branch; // @[Exu.scala 27:19]
  wire  rob_io_branch_info_bits_is_taken; // @[Exu.scala 27:19]
  wire  rob_io_branch_info_bits_predict_miss; // @[Exu.scala 27:19]
  wire  rob_io_need_flush; // @[Exu.scala 27:19]
  wire  alu0_clock; // @[Exu.scala 28:20]
  wire  alu0_reset; // @[Exu.scala 28:20]
  wire  alu0_io_dispatch_info_valid; // @[Exu.scala 28:20]
  wire [5:0] alu0_io_dispatch_info_bits_uop; // @[Exu.scala 28:20]
  wire  alu0_io_dispatch_info_bits_need_imm; // @[Exu.scala 28:20]
  wire [2:0] alu0_io_dispatch_info_bits_rob_idx; // @[Exu.scala 28:20]
  wire [31:0] alu0_io_dispatch_info_bits_op1_data; // @[Exu.scala 28:20]
  wire [31:0] alu0_io_dispatch_info_bits_op2_data; // @[Exu.scala 28:20]
  wire [31:0] alu0_io_dispatch_info_bits_imm_data; // @[Exu.scala 28:20]
  wire  alu0_io_wb_info_valid; // @[Exu.scala 28:20]
  wire [2:0] alu0_io_wb_info_bits_rob_idx; // @[Exu.scala 28:20]
  wire [31:0] alu0_io_wb_info_bits_data; // @[Exu.scala 28:20]
  wire  alu0_io_need_flush; // @[Exu.scala 28:20]
  wire  alu1_clock; // @[Exu.scala 29:20]
  wire  alu1_reset; // @[Exu.scala 29:20]
  wire  alu1_io_dispatch_info_valid; // @[Exu.scala 29:20]
  wire [5:0] alu1_io_dispatch_info_bits_uop; // @[Exu.scala 29:20]
  wire  alu1_io_dispatch_info_bits_need_imm; // @[Exu.scala 29:20]
  wire [2:0] alu1_io_dispatch_info_bits_rob_idx; // @[Exu.scala 29:20]
  wire [31:0] alu1_io_dispatch_info_bits_op1_data; // @[Exu.scala 29:20]
  wire [31:0] alu1_io_dispatch_info_bits_op2_data; // @[Exu.scala 29:20]
  wire [31:0] alu1_io_dispatch_info_bits_imm_data; // @[Exu.scala 29:20]
  wire  alu1_io_wb_info_valid; // @[Exu.scala 29:20]
  wire [2:0] alu1_io_wb_info_bits_rob_idx; // @[Exu.scala 29:20]
  wire [31:0] alu1_io_wb_info_bits_data; // @[Exu.scala 29:20]
  wire  alu1_io_need_flush; // @[Exu.scala 29:20]
  wire  bju0_clock; // @[Exu.scala 31:20]
  wire  bju0_reset; // @[Exu.scala 31:20]
  wire  bju0_io_dispatch_info_valid; // @[Exu.scala 31:20]
  wire [5:0] bju0_io_dispatch_info_bits_uop; // @[Exu.scala 31:20]
  wire [2:0] bju0_io_dispatch_info_bits_rob_idx; // @[Exu.scala 31:20]
  wire [31:0] bju0_io_dispatch_info_bits_inst_addr; // @[Exu.scala 31:20]
  wire [31:0] bju0_io_dispatch_info_bits_op1_data; // @[Exu.scala 31:20]
  wire [31:0] bju0_io_dispatch_info_bits_op2_data; // @[Exu.scala 31:20]
  wire [31:0] bju0_io_dispatch_info_bits_imm_data; // @[Exu.scala 31:20]
  wire  bju0_io_dispatch_info_bits_predict_taken; // @[Exu.scala 31:20]
  wire  bju0_io_wb_info_valid; // @[Exu.scala 31:20]
  wire [2:0] bju0_io_wb_info_bits_rob_idx; // @[Exu.scala 31:20]
  wire [31:0] bju0_io_wb_info_bits_data; // @[Exu.scala 31:20]
  wire [31:0] bju0_io_wb_info_bits_target_addr; // @[Exu.scala 31:20]
  wire  bju0_io_wb_info_bits_is_taken; // @[Exu.scala 31:20]
  wire  bju0_io_wb_info_bits_predict_miss; // @[Exu.scala 31:20]
  wire  bju0_io_need_flush; // @[Exu.scala 31:20]
  wire  lsu_clock; // @[Exu.scala 33:19]
  wire  lsu_reset; // @[Exu.scala 33:19]
  wire  lsu_io_dispatch_info_ready; // @[Exu.scala 33:19]
  wire  lsu_io_dispatch_info_valid; // @[Exu.scala 33:19]
  wire [5:0] lsu_io_dispatch_info_bits_uop; // @[Exu.scala 33:19]
  wire [2:0] lsu_io_dispatch_info_bits_rob_idx; // @[Exu.scala 33:19]
  wire [31:0] lsu_io_dispatch_info_bits_op1_data; // @[Exu.scala 33:19]
  wire [31:0] lsu_io_dispatch_info_bits_op2_data; // @[Exu.scala 33:19]
  wire [31:0] lsu_io_dispatch_info_bits_imm_data; // @[Exu.scala 33:19]
  wire  lsu_io_wb_info_valid; // @[Exu.scala 33:19]
  wire [2:0] lsu_io_wb_info_bits_rob_idx; // @[Exu.scala 33:19]
  wire [31:0] lsu_io_wb_info_bits_data; // @[Exu.scala 33:19]
  wire  lsu_io_rob_commit_0_valid; // @[Exu.scala 33:19]
  wire [2:0] lsu_io_rob_commit_0_bits_des_rob; // @[Exu.scala 33:19]
  wire  lsu_io_rob_commit_1_valid; // @[Exu.scala 33:19]
  wire [2:0] lsu_io_rob_commit_1_bits_des_rob; // @[Exu.scala 33:19]
  wire  lsu_io_cache_read_ready; // @[Exu.scala 33:19]
  wire  lsu_io_cache_read_valid; // @[Exu.scala 33:19]
  wire [31:0] lsu_io_cache_read_bits_addr; // @[Exu.scala 33:19]
  wire [3:0] lsu_io_cache_read_bits_rob_idx; // @[Exu.scala 33:19]
  wire  lsu_io_cache_write_ready; // @[Exu.scala 33:19]
  wire  lsu_io_cache_write_valid; // @[Exu.scala 33:19]
  wire [31:0] lsu_io_cache_write_bits_addr; // @[Exu.scala 33:19]
  wire [31:0] lsu_io_cache_write_bits_data; // @[Exu.scala 33:19]
  wire [3:0] lsu_io_cache_write_bits_byte_mask; // @[Exu.scala 33:19]
  wire [31:0] lsu_io_cache_resp_data; // @[Exu.scala 33:19]
  wire  lsu_io_need_flush; // @[Exu.scala 33:19]
  wire  mdu_clock; // @[Exu.scala 34:19]
  wire  mdu_reset; // @[Exu.scala 34:19]
  wire  mdu_io_dispatch_info_valid; // @[Exu.scala 34:19]
  wire [2:0] mdu_io_dispatch_info_bits_rob_idx; // @[Exu.scala 34:19]
  wire [31:0] mdu_io_dispatch_info_bits_op1_data; // @[Exu.scala 34:19]
  wire [31:0] mdu_io_dispatch_info_bits_op2_data; // @[Exu.scala 34:19]
  wire  mdu_io_wb_info_valid; // @[Exu.scala 34:19]
  wire [2:0] mdu_io_wb_info_bits_rob_idx; // @[Exu.scala 34:19]
  wire [31:0] mdu_io_wb_info_bits_data; // @[Exu.scala 34:19]
  wire  mdu_io_need_flush; // @[Exu.scala 34:19]
  wire  dcache_io_dcache_read_req_ready; // @[Exu.scala 35:22]
  wire  dcache_io_dcache_read_req_valid; // @[Exu.scala 35:22]
  wire [31:0] dcache_io_dcache_read_req_bits_addr; // @[Exu.scala 35:22]
  wire [3:0] dcache_io_dcache_read_req_bits_rob_idx; // @[Exu.scala 35:22]
  wire [31:0] dcache_io_dcache_read_resp_data; // @[Exu.scala 35:22]
  wire  dcache_io_dcache_write_req_ready; // @[Exu.scala 35:22]
  wire  dcache_io_dcache_write_req_valid; // @[Exu.scala 35:22]
  wire [31:0] dcache_io_dcache_write_req_bits_addr; // @[Exu.scala 35:22]
  wire [31:0] dcache_io_dcache_write_req_bits_data; // @[Exu.scala 35:22]
  wire [3:0] dcache_io_dcache_write_req_bits_byte_mask; // @[Exu.scala 35:22]
  wire  dcache_io_io_read_req_ready; // @[Exu.scala 35:22]
  wire  dcache_io_io_read_req_valid; // @[Exu.scala 35:22]
  wire [31:0] dcache_io_io_read_req_bits_addr; // @[Exu.scala 35:22]
  wire [3:0] dcache_io_io_read_req_bits_rob_idx; // @[Exu.scala 35:22]
  wire [31:0] dcache_io_io_read_resp_bits_data; // @[Exu.scala 35:22]
  wire  dcache_io_io_write_req_ready; // @[Exu.scala 35:22]
  wire  dcache_io_io_write_req_valid; // @[Exu.scala 35:22]
  wire [31:0] dcache_io_io_write_req_bits_addr; // @[Exu.scala 35:22]
  wire [31:0] dcache_io_io_write_req_bits_data; // @[Exu.scala 35:22]
  wire [3:0] dcache_io_io_write_req_bits_byte_mask; // @[Exu.scala 35:22]
  Decode decode ( // @[Exu.scala 24:22]
    .clock(decode_clock),
    .reset(decode_reset),
    .io_fb_inst_bank_valid(decode_io_fb_inst_bank_valid),
    .io_fb_inst_bank_bits_data_0_inst(decode_io_fb_inst_bank_bits_data_0_inst),
    .io_fb_inst_bank_bits_data_0_inst_addr(decode_io_fb_inst_bank_bits_data_0_inst_addr),
    .io_fb_inst_bank_bits_data_0_gh_backup(decode_io_fb_inst_bank_bits_data_0_gh_backup),
    .io_fb_inst_bank_bits_data_0_is_valid(decode_io_fb_inst_bank_bits_data_0_is_valid),
    .io_fb_inst_bank_bits_data_0_predict_taken(decode_io_fb_inst_bank_bits_data_0_predict_taken),
    .io_fb_inst_bank_bits_data_1_inst(decode_io_fb_inst_bank_bits_data_1_inst),
    .io_fb_inst_bank_bits_data_1_inst_addr(decode_io_fb_inst_bank_bits_data_1_inst_addr),
    .io_fb_inst_bank_bits_data_1_gh_backup(decode_io_fb_inst_bank_bits_data_1_gh_backup),
    .io_fb_inst_bank_bits_data_1_is_valid(decode_io_fb_inst_bank_bits_data_1_is_valid),
    .io_fb_inst_bank_bits_data_1_predict_taken(decode_io_fb_inst_bank_bits_data_1_predict_taken),
    .io_fb_resp_deq_valid_0(decode_io_fb_resp_deq_valid_0),
    .io_fb_resp_deq_valid_1(decode_io_fb_resp_deq_valid_1),
    .io_rob_allocate_allocate_req_valid(decode_io_rob_allocate_allocate_req_valid),
    .io_rob_allocate_allocate_req_bits_0(decode_io_rob_allocate_allocate_req_bits_0),
    .io_rob_allocate_allocate_req_bits_1(decode_io_rob_allocate_allocate_req_bits_1),
    .io_rob_allocate_allocate_info_valid(decode_io_rob_allocate_allocate_info_valid),
    .io_rob_allocate_allocate_info_bits_0_rob_idx(decode_io_rob_allocate_allocate_info_bits_0_rob_idx),
    .io_rob_allocate_allocate_info_bits_0_inst_valid(decode_io_rob_allocate_allocate_info_bits_0_inst_valid),
    .io_rob_allocate_allocate_info_bits_0_inst_addr(decode_io_rob_allocate_allocate_info_bits_0_inst_addr),
    .io_rob_allocate_allocate_info_bits_0_uop(decode_io_rob_allocate_allocate_info_bits_0_uop),
    .io_rob_allocate_allocate_info_bits_0_unit_sel(decode_io_rob_allocate_allocate_info_bits_0_unit_sel),
    .io_rob_allocate_allocate_info_bits_0_need_imm(decode_io_rob_allocate_allocate_info_bits_0_need_imm),
    .io_rob_allocate_allocate_info_bits_0_commit_addr(decode_io_rob_allocate_allocate_info_bits_0_commit_addr),
    .io_rob_allocate_allocate_info_bits_0_gh_info(decode_io_rob_allocate_allocate_info_bits_0_gh_info),
    .io_rob_allocate_allocate_info_bits_0_imm_data(decode_io_rob_allocate_allocate_info_bits_0_imm_data),
    .io_rob_allocate_allocate_info_bits_0_flush_on_commit(decode_io_rob_allocate_allocate_info_bits_0_flush_on_commit),
    .io_rob_allocate_allocate_info_bits_0_predict_taken(decode_io_rob_allocate_allocate_info_bits_0_predict_taken),
    .io_rob_allocate_allocate_info_bits_1_rob_idx(decode_io_rob_allocate_allocate_info_bits_1_rob_idx),
    .io_rob_allocate_allocate_info_bits_1_inst_valid(decode_io_rob_allocate_allocate_info_bits_1_inst_valid),
    .io_rob_allocate_allocate_info_bits_1_inst_addr(decode_io_rob_allocate_allocate_info_bits_1_inst_addr),
    .io_rob_allocate_allocate_info_bits_1_uop(decode_io_rob_allocate_allocate_info_bits_1_uop),
    .io_rob_allocate_allocate_info_bits_1_unit_sel(decode_io_rob_allocate_allocate_info_bits_1_unit_sel),
    .io_rob_allocate_allocate_info_bits_1_need_imm(decode_io_rob_allocate_allocate_info_bits_1_need_imm),
    .io_rob_allocate_allocate_info_bits_1_commit_addr(decode_io_rob_allocate_allocate_info_bits_1_commit_addr),
    .io_rob_allocate_allocate_info_bits_1_gh_info(decode_io_rob_allocate_allocate_info_bits_1_gh_info),
    .io_rob_allocate_allocate_info_bits_1_imm_data(decode_io_rob_allocate_allocate_info_bits_1_imm_data),
    .io_rob_allocate_allocate_info_bits_1_flush_on_commit(decode_io_rob_allocate_allocate_info_bits_1_flush_on_commit),
    .io_rob_allocate_allocate_info_bits_1_predict_taken(decode_io_rob_allocate_allocate_info_bits_1_predict_taken),
    .io_rob_allocate_allocate_resp_valid(decode_io_rob_allocate_allocate_resp_valid),
    .io_rob_allocate_allocate_resp_bits_rob_idx_0(decode_io_rob_allocate_allocate_resp_bits_rob_idx_0),
    .io_rob_allocate_allocate_resp_bits_rob_idx_1(decode_io_rob_allocate_allocate_resp_bits_rob_idx_1),
    .io_rob_allocate_allocate_resp_bits_enq_valid_mask_0(decode_io_rob_allocate_allocate_resp_bits_enq_valid_mask_0),
    .io_rob_allocate_allocate_resp_bits_enq_valid_mask_1(decode_io_rob_allocate_allocate_resp_bits_enq_valid_mask_1),
    .io_rename_info_valid(decode_io_rename_info_valid),
    .io_rename_info_bits_0_is_valid(decode_io_rename_info_bits_0_is_valid),
    .io_rename_info_bits_0_op1_addr(decode_io_rename_info_bits_0_op1_addr),
    .io_rename_info_bits_0_op2_addr(decode_io_rename_info_bits_0_op2_addr),
    .io_rename_info_bits_0_des_addr(decode_io_rename_info_bits_0_des_addr),
    .io_rename_info_bits_0_des_rob(decode_io_rename_info_bits_0_des_rob),
    .io_rename_info_bits_1_is_valid(decode_io_rename_info_bits_1_is_valid),
    .io_rename_info_bits_1_op1_addr(decode_io_rename_info_bits_1_op1_addr),
    .io_rename_info_bits_1_op2_addr(decode_io_rename_info_bits_1_op2_addr),
    .io_rename_info_bits_1_des_addr(decode_io_rename_info_bits_1_des_addr),
    .io_rename_info_bits_1_des_rob(decode_io_rename_info_bits_1_des_rob),
    .io_need_flush(decode_io_need_flush)
  );
  Rename rename ( // @[Exu.scala 25:22]
    .clock(rename_clock),
    .reset(rename_reset),
    .io_rename_info_valid(rename_io_rename_info_valid),
    .io_rename_info_bits_0_is_valid(rename_io_rename_info_bits_0_is_valid),
    .io_rename_info_bits_0_op1_addr(rename_io_rename_info_bits_0_op1_addr),
    .io_rename_info_bits_0_op2_addr(rename_io_rename_info_bits_0_op2_addr),
    .io_rename_info_bits_0_des_addr(rename_io_rename_info_bits_0_des_addr),
    .io_rename_info_bits_0_des_rob(rename_io_rename_info_bits_0_des_rob),
    .io_rename_info_bits_1_is_valid(rename_io_rename_info_bits_1_is_valid),
    .io_rename_info_bits_1_op1_addr(rename_io_rename_info_bits_1_op1_addr),
    .io_rename_info_bits_1_op2_addr(rename_io_rename_info_bits_1_op2_addr),
    .io_rename_info_bits_1_des_addr(rename_io_rename_info_bits_1_des_addr),
    .io_rename_info_bits_1_des_rob(rename_io_rename_info_bits_1_des_rob),
    .io_rob_commit_0_valid(rename_io_rob_commit_0_valid),
    .io_rob_commit_0_bits_des_rob(rename_io_rob_commit_0_bits_des_rob),
    .io_rob_commit_0_bits_commit_addr(rename_io_rob_commit_0_bits_commit_addr),
    .io_rob_commit_1_valid(rename_io_rob_commit_1_valid),
    .io_rob_commit_1_bits_des_rob(rename_io_rob_commit_1_bits_des_rob),
    .io_rob_commit_1_bits_commit_addr(rename_io_rob_commit_1_bits_commit_addr),
    .io_reg_read_0_op1_addr(rename_io_reg_read_0_op1_addr),
    .io_reg_read_0_op2_addr(rename_io_reg_read_0_op2_addr),
    .io_reg_read_0_op1_data(rename_io_reg_read_0_op1_data),
    .io_reg_read_0_op2_data(rename_io_reg_read_0_op2_data),
    .io_reg_read_1_op1_addr(rename_io_reg_read_1_op1_addr),
    .io_reg_read_1_op2_addr(rename_io_reg_read_1_op2_addr),
    .io_reg_read_1_op1_data(rename_io_reg_read_1_op1_data),
    .io_reg_read_1_op2_data(rename_io_reg_read_1_op2_data),
    .io_rob_init_info_valid(rename_io_rob_init_info_valid),
    .io_rob_init_info_bits_0_is_valid(rename_io_rob_init_info_bits_0_is_valid),
    .io_rob_init_info_bits_0_des_rob(rename_io_rob_init_info_bits_0_des_rob),
    .io_rob_init_info_bits_0_op1_rob(rename_io_rob_init_info_bits_0_op1_rob),
    .io_rob_init_info_bits_0_op2_rob(rename_io_rob_init_info_bits_0_op2_rob),
    .io_rob_init_info_bits_0_op1_regData(rename_io_rob_init_info_bits_0_op1_regData),
    .io_rob_init_info_bits_0_op2_regData(rename_io_rob_init_info_bits_0_op2_regData),
    .io_rob_init_info_bits_0_op1_in_rob(rename_io_rob_init_info_bits_0_op1_in_rob),
    .io_rob_init_info_bits_0_op2_in_rob(rename_io_rob_init_info_bits_0_op2_in_rob),
    .io_rob_init_info_bits_1_is_valid(rename_io_rob_init_info_bits_1_is_valid),
    .io_rob_init_info_bits_1_des_rob(rename_io_rob_init_info_bits_1_des_rob),
    .io_rob_init_info_bits_1_op1_rob(rename_io_rob_init_info_bits_1_op1_rob),
    .io_rob_init_info_bits_1_op2_rob(rename_io_rob_init_info_bits_1_op2_rob),
    .io_rob_init_info_bits_1_op1_regData(rename_io_rob_init_info_bits_1_op1_regData),
    .io_rob_init_info_bits_1_op2_regData(rename_io_rob_init_info_bits_1_op2_regData),
    .io_rob_init_info_bits_1_op1_in_rob(rename_io_rob_init_info_bits_1_op1_in_rob),
    .io_rob_init_info_bits_1_op2_in_rob(rename_io_rob_init_info_bits_1_op2_in_rob),
    .io_need_flush(rename_io_need_flush)
  );
  Regfile regfile ( // @[Exu.scala 26:23]
    .clock(regfile_clock),
    .reset(regfile_reset),
    .io_reg_read_0_op1_addr(regfile_io_reg_read_0_op1_addr),
    .io_reg_read_0_op2_addr(regfile_io_reg_read_0_op2_addr),
    .io_reg_read_0_op1_data(regfile_io_reg_read_0_op1_data),
    .io_reg_read_0_op2_data(regfile_io_reg_read_0_op2_data),
    .io_reg_read_1_op1_addr(regfile_io_reg_read_1_op1_addr),
    .io_reg_read_1_op2_addr(regfile_io_reg_read_1_op2_addr),
    .io_reg_read_1_op1_data(regfile_io_reg_read_1_op1_data),
    .io_reg_read_1_op2_data(regfile_io_reg_read_1_op2_data),
    .io_rob_commit_i_0_valid(regfile_io_rob_commit_i_0_valid),
    .io_rob_commit_i_0_bits_commit_addr(regfile_io_rob_commit_i_0_bits_commit_addr),
    .io_rob_commit_i_0_bits_commit_data(regfile_io_rob_commit_i_0_bits_commit_data),
    .io_rob_commit_i_1_valid(regfile_io_rob_commit_i_1_valid),
    .io_rob_commit_i_1_bits_commit_addr(regfile_io_rob_commit_i_1_bits_commit_addr),
    .io_rob_commit_i_1_bits_commit_data(regfile_io_rob_commit_i_1_bits_commit_data)
  );
  Rob rob ( // @[Exu.scala 27:19]
    .clock(rob_clock),
    .reset(rob_reset),
    .io_rob_allocate_allocate_req_valid(rob_io_rob_allocate_allocate_req_valid),
    .io_rob_allocate_allocate_req_bits_0(rob_io_rob_allocate_allocate_req_bits_0),
    .io_rob_allocate_allocate_req_bits_1(rob_io_rob_allocate_allocate_req_bits_1),
    .io_rob_allocate_allocate_info_valid(rob_io_rob_allocate_allocate_info_valid),
    .io_rob_allocate_allocate_info_bits_0_rob_idx(rob_io_rob_allocate_allocate_info_bits_0_rob_idx),
    .io_rob_allocate_allocate_info_bits_0_inst_valid(rob_io_rob_allocate_allocate_info_bits_0_inst_valid),
    .io_rob_allocate_allocate_info_bits_0_inst_addr(rob_io_rob_allocate_allocate_info_bits_0_inst_addr),
    .io_rob_allocate_allocate_info_bits_0_uop(rob_io_rob_allocate_allocate_info_bits_0_uop),
    .io_rob_allocate_allocate_info_bits_0_unit_sel(rob_io_rob_allocate_allocate_info_bits_0_unit_sel),
    .io_rob_allocate_allocate_info_bits_0_need_imm(rob_io_rob_allocate_allocate_info_bits_0_need_imm),
    .io_rob_allocate_allocate_info_bits_0_commit_addr(rob_io_rob_allocate_allocate_info_bits_0_commit_addr),
    .io_rob_allocate_allocate_info_bits_0_gh_info(rob_io_rob_allocate_allocate_info_bits_0_gh_info),
    .io_rob_allocate_allocate_info_bits_0_imm_data(rob_io_rob_allocate_allocate_info_bits_0_imm_data),
    .io_rob_allocate_allocate_info_bits_0_flush_on_commit(rob_io_rob_allocate_allocate_info_bits_0_flush_on_commit),
    .io_rob_allocate_allocate_info_bits_0_predict_taken(rob_io_rob_allocate_allocate_info_bits_0_predict_taken),
    .io_rob_allocate_allocate_info_bits_1_rob_idx(rob_io_rob_allocate_allocate_info_bits_1_rob_idx),
    .io_rob_allocate_allocate_info_bits_1_inst_valid(rob_io_rob_allocate_allocate_info_bits_1_inst_valid),
    .io_rob_allocate_allocate_info_bits_1_inst_addr(rob_io_rob_allocate_allocate_info_bits_1_inst_addr),
    .io_rob_allocate_allocate_info_bits_1_uop(rob_io_rob_allocate_allocate_info_bits_1_uop),
    .io_rob_allocate_allocate_info_bits_1_unit_sel(rob_io_rob_allocate_allocate_info_bits_1_unit_sel),
    .io_rob_allocate_allocate_info_bits_1_need_imm(rob_io_rob_allocate_allocate_info_bits_1_need_imm),
    .io_rob_allocate_allocate_info_bits_1_commit_addr(rob_io_rob_allocate_allocate_info_bits_1_commit_addr),
    .io_rob_allocate_allocate_info_bits_1_gh_info(rob_io_rob_allocate_allocate_info_bits_1_gh_info),
    .io_rob_allocate_allocate_info_bits_1_imm_data(rob_io_rob_allocate_allocate_info_bits_1_imm_data),
    .io_rob_allocate_allocate_info_bits_1_flush_on_commit(rob_io_rob_allocate_allocate_info_bits_1_flush_on_commit),
    .io_rob_allocate_allocate_info_bits_1_predict_taken(rob_io_rob_allocate_allocate_info_bits_1_predict_taken),
    .io_rob_allocate_allocate_resp_valid(rob_io_rob_allocate_allocate_resp_valid),
    .io_rob_allocate_allocate_resp_bits_rob_idx_0(rob_io_rob_allocate_allocate_resp_bits_rob_idx_0),
    .io_rob_allocate_allocate_resp_bits_rob_idx_1(rob_io_rob_allocate_allocate_resp_bits_rob_idx_1),
    .io_rob_allocate_allocate_resp_bits_enq_valid_mask_0(rob_io_rob_allocate_allocate_resp_bits_enq_valid_mask_0),
    .io_rob_allocate_allocate_resp_bits_enq_valid_mask_1(rob_io_rob_allocate_allocate_resp_bits_enq_valid_mask_1),
    .io_rob_init_info_valid(rob_io_rob_init_info_valid),
    .io_rob_init_info_bits_0_is_valid(rob_io_rob_init_info_bits_0_is_valid),
    .io_rob_init_info_bits_0_des_rob(rob_io_rob_init_info_bits_0_des_rob),
    .io_rob_init_info_bits_0_op1_rob(rob_io_rob_init_info_bits_0_op1_rob),
    .io_rob_init_info_bits_0_op2_rob(rob_io_rob_init_info_bits_0_op2_rob),
    .io_rob_init_info_bits_0_op1_regData(rob_io_rob_init_info_bits_0_op1_regData),
    .io_rob_init_info_bits_0_op2_regData(rob_io_rob_init_info_bits_0_op2_regData),
    .io_rob_init_info_bits_0_op1_in_rob(rob_io_rob_init_info_bits_0_op1_in_rob),
    .io_rob_init_info_bits_0_op2_in_rob(rob_io_rob_init_info_bits_0_op2_in_rob),
    .io_rob_init_info_bits_1_is_valid(rob_io_rob_init_info_bits_1_is_valid),
    .io_rob_init_info_bits_1_des_rob(rob_io_rob_init_info_bits_1_des_rob),
    .io_rob_init_info_bits_1_op1_rob(rob_io_rob_init_info_bits_1_op1_rob),
    .io_rob_init_info_bits_1_op2_rob(rob_io_rob_init_info_bits_1_op2_rob),
    .io_rob_init_info_bits_1_op1_regData(rob_io_rob_init_info_bits_1_op1_regData),
    .io_rob_init_info_bits_1_op2_regData(rob_io_rob_init_info_bits_1_op2_regData),
    .io_rob_init_info_bits_1_op1_in_rob(rob_io_rob_init_info_bits_1_op1_in_rob),
    .io_rob_init_info_bits_1_op2_in_rob(rob_io_rob_init_info_bits_1_op2_in_rob),
    .io_wb_info_i_0_valid(rob_io_wb_info_i_0_valid),
    .io_wb_info_i_0_bits_rob_idx(rob_io_wb_info_i_0_bits_rob_idx),
    .io_wb_info_i_0_bits_data(rob_io_wb_info_i_0_bits_data),
    .io_wb_info_i_1_valid(rob_io_wb_info_i_1_valid),
    .io_wb_info_i_1_bits_rob_idx(rob_io_wb_info_i_1_bits_rob_idx),
    .io_wb_info_i_1_bits_data(rob_io_wb_info_i_1_bits_data),
    .io_wb_info_i_2_valid(rob_io_wb_info_i_2_valid),
    .io_wb_info_i_2_bits_rob_idx(rob_io_wb_info_i_2_bits_rob_idx),
    .io_wb_info_i_2_bits_data(rob_io_wb_info_i_2_bits_data),
    .io_wb_info_i_2_bits_target_addr(rob_io_wb_info_i_2_bits_target_addr),
    .io_wb_info_i_2_bits_is_taken(rob_io_wb_info_i_2_bits_is_taken),
    .io_wb_info_i_2_bits_predict_miss(rob_io_wb_info_i_2_bits_predict_miss),
    .io_wb_info_i_3_valid(rob_io_wb_info_i_3_valid),
    .io_wb_info_i_3_bits_rob_idx(rob_io_wb_info_i_3_bits_rob_idx),
    .io_wb_info_i_3_bits_data(rob_io_wb_info_i_3_bits_data),
    .io_wb_info_i_4_valid(rob_io_wb_info_i_4_valid),
    .io_wb_info_i_4_bits_rob_idx(rob_io_wb_info_i_4_bits_rob_idx),
    .io_wb_info_i_4_bits_data(rob_io_wb_info_i_4_bits_data),
    .io_dispatch_info_o_0_valid(rob_io_dispatch_info_o_0_valid),
    .io_dispatch_info_o_0_bits_uop(rob_io_dispatch_info_o_0_bits_uop),
    .io_dispatch_info_o_0_bits_need_imm(rob_io_dispatch_info_o_0_bits_need_imm),
    .io_dispatch_info_o_0_bits_rob_idx(rob_io_dispatch_info_o_0_bits_rob_idx),
    .io_dispatch_info_o_0_bits_op1_data(rob_io_dispatch_info_o_0_bits_op1_data),
    .io_dispatch_info_o_0_bits_op2_data(rob_io_dispatch_info_o_0_bits_op2_data),
    .io_dispatch_info_o_0_bits_imm_data(rob_io_dispatch_info_o_0_bits_imm_data),
    .io_dispatch_info_o_1_valid(rob_io_dispatch_info_o_1_valid),
    .io_dispatch_info_o_1_bits_uop(rob_io_dispatch_info_o_1_bits_uop),
    .io_dispatch_info_o_1_bits_need_imm(rob_io_dispatch_info_o_1_bits_need_imm),
    .io_dispatch_info_o_1_bits_rob_idx(rob_io_dispatch_info_o_1_bits_rob_idx),
    .io_dispatch_info_o_1_bits_op1_data(rob_io_dispatch_info_o_1_bits_op1_data),
    .io_dispatch_info_o_1_bits_op2_data(rob_io_dispatch_info_o_1_bits_op2_data),
    .io_dispatch_info_o_1_bits_imm_data(rob_io_dispatch_info_o_1_bits_imm_data),
    .io_dispatch_info_o_2_valid(rob_io_dispatch_info_o_2_valid),
    .io_dispatch_info_o_2_bits_uop(rob_io_dispatch_info_o_2_bits_uop),
    .io_dispatch_info_o_2_bits_rob_idx(rob_io_dispatch_info_o_2_bits_rob_idx),
    .io_dispatch_info_o_2_bits_inst_addr(rob_io_dispatch_info_o_2_bits_inst_addr),
    .io_dispatch_info_o_2_bits_op1_data(rob_io_dispatch_info_o_2_bits_op1_data),
    .io_dispatch_info_o_2_bits_op2_data(rob_io_dispatch_info_o_2_bits_op2_data),
    .io_dispatch_info_o_2_bits_imm_data(rob_io_dispatch_info_o_2_bits_imm_data),
    .io_dispatch_info_o_2_bits_predict_taken(rob_io_dispatch_info_o_2_bits_predict_taken),
    .io_dispatch_info_o_3_valid(rob_io_dispatch_info_o_3_valid),
    .io_dispatch_info_o_3_bits_rob_idx(rob_io_dispatch_info_o_3_bits_rob_idx),
    .io_dispatch_info_o_3_bits_op1_data(rob_io_dispatch_info_o_3_bits_op1_data),
    .io_dispatch_info_o_3_bits_op2_data(rob_io_dispatch_info_o_3_bits_op2_data),
    .io_dispatch_info_o_4_ready(rob_io_dispatch_info_o_4_ready),
    .io_dispatch_info_o_4_valid(rob_io_dispatch_info_o_4_valid),
    .io_dispatch_info_o_4_bits_uop(rob_io_dispatch_info_o_4_bits_uop),
    .io_dispatch_info_o_4_bits_rob_idx(rob_io_dispatch_info_o_4_bits_rob_idx),
    .io_dispatch_info_o_4_bits_op1_data(rob_io_dispatch_info_o_4_bits_op1_data),
    .io_dispatch_info_o_4_bits_op2_data(rob_io_dispatch_info_o_4_bits_op2_data),
    .io_dispatch_info_o_4_bits_imm_data(rob_io_dispatch_info_o_4_bits_imm_data),
    .io_rob_commit_0_valid(rob_io_rob_commit_0_valid),
    .io_rob_commit_0_bits_des_rob(rob_io_rob_commit_0_bits_des_rob),
    .io_rob_commit_0_bits_commit_addr(rob_io_rob_commit_0_bits_commit_addr),
    .io_rob_commit_0_bits_commit_data(rob_io_rob_commit_0_bits_commit_data),
    .io_rob_commit_1_valid(rob_io_rob_commit_1_valid),
    .io_rob_commit_1_bits_des_rob(rob_io_rob_commit_1_bits_des_rob),
    .io_rob_commit_1_bits_commit_addr(rob_io_rob_commit_1_bits_commit_addr),
    .io_rob_commit_1_bits_commit_data(rob_io_rob_commit_1_bits_commit_data),
    .io_branch_info_valid(rob_io_branch_info_valid),
    .io_branch_info_bits_target_addr(rob_io_branch_info_bits_target_addr),
    .io_branch_info_bits_inst_addr(rob_io_branch_info_bits_inst_addr),
    .io_branch_info_bits_gh_update(rob_io_branch_info_bits_gh_update),
    .io_branch_info_bits_is_branch(rob_io_branch_info_bits_is_branch),
    .io_branch_info_bits_is_taken(rob_io_branch_info_bits_is_taken),
    .io_branch_info_bits_predict_miss(rob_io_branch_info_bits_predict_miss),
    .io_need_flush(rob_io_need_flush)
  );
  Alu alu0 ( // @[Exu.scala 28:20]
    .clock(alu0_clock),
    .reset(alu0_reset),
    .io_dispatch_info_valid(alu0_io_dispatch_info_valid),
    .io_dispatch_info_bits_uop(alu0_io_dispatch_info_bits_uop),
    .io_dispatch_info_bits_need_imm(alu0_io_dispatch_info_bits_need_imm),
    .io_dispatch_info_bits_rob_idx(alu0_io_dispatch_info_bits_rob_idx),
    .io_dispatch_info_bits_op1_data(alu0_io_dispatch_info_bits_op1_data),
    .io_dispatch_info_bits_op2_data(alu0_io_dispatch_info_bits_op2_data),
    .io_dispatch_info_bits_imm_data(alu0_io_dispatch_info_bits_imm_data),
    .io_wb_info_valid(alu0_io_wb_info_valid),
    .io_wb_info_bits_rob_idx(alu0_io_wb_info_bits_rob_idx),
    .io_wb_info_bits_data(alu0_io_wb_info_bits_data),
    .io_need_flush(alu0_io_need_flush)
  );
  Alu alu1 ( // @[Exu.scala 29:20]
    .clock(alu1_clock),
    .reset(alu1_reset),
    .io_dispatch_info_valid(alu1_io_dispatch_info_valid),
    .io_dispatch_info_bits_uop(alu1_io_dispatch_info_bits_uop),
    .io_dispatch_info_bits_need_imm(alu1_io_dispatch_info_bits_need_imm),
    .io_dispatch_info_bits_rob_idx(alu1_io_dispatch_info_bits_rob_idx),
    .io_dispatch_info_bits_op1_data(alu1_io_dispatch_info_bits_op1_data),
    .io_dispatch_info_bits_op2_data(alu1_io_dispatch_info_bits_op2_data),
    .io_dispatch_info_bits_imm_data(alu1_io_dispatch_info_bits_imm_data),
    .io_wb_info_valid(alu1_io_wb_info_valid),
    .io_wb_info_bits_rob_idx(alu1_io_wb_info_bits_rob_idx),
    .io_wb_info_bits_data(alu1_io_wb_info_bits_data),
    .io_need_flush(alu1_io_need_flush)
  );
  Bju bju0 ( // @[Exu.scala 31:20]
    .clock(bju0_clock),
    .reset(bju0_reset),
    .io_dispatch_info_valid(bju0_io_dispatch_info_valid),
    .io_dispatch_info_bits_uop(bju0_io_dispatch_info_bits_uop),
    .io_dispatch_info_bits_rob_idx(bju0_io_dispatch_info_bits_rob_idx),
    .io_dispatch_info_bits_inst_addr(bju0_io_dispatch_info_bits_inst_addr),
    .io_dispatch_info_bits_op1_data(bju0_io_dispatch_info_bits_op1_data),
    .io_dispatch_info_bits_op2_data(bju0_io_dispatch_info_bits_op2_data),
    .io_dispatch_info_bits_imm_data(bju0_io_dispatch_info_bits_imm_data),
    .io_dispatch_info_bits_predict_taken(bju0_io_dispatch_info_bits_predict_taken),
    .io_wb_info_valid(bju0_io_wb_info_valid),
    .io_wb_info_bits_rob_idx(bju0_io_wb_info_bits_rob_idx),
    .io_wb_info_bits_data(bju0_io_wb_info_bits_data),
    .io_wb_info_bits_target_addr(bju0_io_wb_info_bits_target_addr),
    .io_wb_info_bits_is_taken(bju0_io_wb_info_bits_is_taken),
    .io_wb_info_bits_predict_miss(bju0_io_wb_info_bits_predict_miss),
    .io_need_flush(bju0_io_need_flush)
  );
  Lsu lsu ( // @[Exu.scala 33:19]
    .clock(lsu_clock),
    .reset(lsu_reset),
    .io_dispatch_info_ready(lsu_io_dispatch_info_ready),
    .io_dispatch_info_valid(lsu_io_dispatch_info_valid),
    .io_dispatch_info_bits_uop(lsu_io_dispatch_info_bits_uop),
    .io_dispatch_info_bits_rob_idx(lsu_io_dispatch_info_bits_rob_idx),
    .io_dispatch_info_bits_op1_data(lsu_io_dispatch_info_bits_op1_data),
    .io_dispatch_info_bits_op2_data(lsu_io_dispatch_info_bits_op2_data),
    .io_dispatch_info_bits_imm_data(lsu_io_dispatch_info_bits_imm_data),
    .io_wb_info_valid(lsu_io_wb_info_valid),
    .io_wb_info_bits_rob_idx(lsu_io_wb_info_bits_rob_idx),
    .io_wb_info_bits_data(lsu_io_wb_info_bits_data),
    .io_rob_commit_0_valid(lsu_io_rob_commit_0_valid),
    .io_rob_commit_0_bits_des_rob(lsu_io_rob_commit_0_bits_des_rob),
    .io_rob_commit_1_valid(lsu_io_rob_commit_1_valid),
    .io_rob_commit_1_bits_des_rob(lsu_io_rob_commit_1_bits_des_rob),
    .io_cache_read_ready(lsu_io_cache_read_ready),
    .io_cache_read_valid(lsu_io_cache_read_valid),
    .io_cache_read_bits_addr(lsu_io_cache_read_bits_addr),
    .io_cache_read_bits_rob_idx(lsu_io_cache_read_bits_rob_idx),
    .io_cache_write_ready(lsu_io_cache_write_ready),
    .io_cache_write_valid(lsu_io_cache_write_valid),
    .io_cache_write_bits_addr(lsu_io_cache_write_bits_addr),
    .io_cache_write_bits_data(lsu_io_cache_write_bits_data),
    .io_cache_write_bits_byte_mask(lsu_io_cache_write_bits_byte_mask),
    .io_cache_resp_data(lsu_io_cache_resp_data),
    .io_need_flush(lsu_io_need_flush)
  );
  Mdu mdu ( // @[Exu.scala 34:19]
    .clock(mdu_clock),
    .reset(mdu_reset),
    .io_dispatch_info_valid(mdu_io_dispatch_info_valid),
    .io_dispatch_info_bits_rob_idx(mdu_io_dispatch_info_bits_rob_idx),
    .io_dispatch_info_bits_op1_data(mdu_io_dispatch_info_bits_op1_data),
    .io_dispatch_info_bits_op2_data(mdu_io_dispatch_info_bits_op2_data),
    .io_wb_info_valid(mdu_io_wb_info_valid),
    .io_wb_info_bits_rob_idx(mdu_io_wb_info_bits_rob_idx),
    .io_wb_info_bits_data(mdu_io_wb_info_bits_data),
    .io_need_flush(mdu_io_need_flush)
  );
  Dcache dcache ( // @[Exu.scala 35:22]
    .io_dcache_read_req_ready(dcache_io_dcache_read_req_ready),
    .io_dcache_read_req_valid(dcache_io_dcache_read_req_valid),
    .io_dcache_read_req_bits_addr(dcache_io_dcache_read_req_bits_addr),
    .io_dcache_read_req_bits_rob_idx(dcache_io_dcache_read_req_bits_rob_idx),
    .io_dcache_read_resp_data(dcache_io_dcache_read_resp_data),
    .io_dcache_write_req_ready(dcache_io_dcache_write_req_ready),
    .io_dcache_write_req_valid(dcache_io_dcache_write_req_valid),
    .io_dcache_write_req_bits_addr(dcache_io_dcache_write_req_bits_addr),
    .io_dcache_write_req_bits_data(dcache_io_dcache_write_req_bits_data),
    .io_dcache_write_req_bits_byte_mask(dcache_io_dcache_write_req_bits_byte_mask),
    .io_io_read_req_ready(dcache_io_io_read_req_ready),
    .io_io_read_req_valid(dcache_io_io_read_req_valid),
    .io_io_read_req_bits_addr(dcache_io_io_read_req_bits_addr),
    .io_io_read_req_bits_rob_idx(dcache_io_io_read_req_bits_rob_idx),
    .io_io_read_resp_bits_data(dcache_io_io_read_resp_bits_data),
    .io_io_write_req_ready(dcache_io_io_write_req_ready),
    .io_io_write_req_valid(dcache_io_io_write_req_valid),
    .io_io_write_req_bits_addr(dcache_io_io_write_req_bits_addr),
    .io_io_write_req_bits_data(dcache_io_io_write_req_bits_data),
    .io_io_write_req_bits_byte_mask(dcache_io_io_write_req_bits_byte_mask)
  );
  assign io_fb_resp_deq_valid_0 = decode_io_fb_resp_deq_valid_0; // @[Exu.scala 38:20]
  assign io_fb_resp_deq_valid_1 = decode_io_fb_resp_deq_valid_1; // @[Exu.scala 38:20]
  assign io_ex_branch_info_o_valid = rob_io_branch_info_valid; // @[Exu.scala 46:22]
  assign io_ex_branch_info_o_bits_target_addr = rob_io_branch_info_bits_target_addr; // @[Exu.scala 46:22]
  assign io_ex_branch_info_o_bits_inst_addr = rob_io_branch_info_bits_inst_addr; // @[Exu.scala 46:22]
  assign io_ex_branch_info_o_bits_gh_update = rob_io_branch_info_bits_gh_update; // @[Exu.scala 46:22]
  assign io_ex_branch_info_o_bits_is_branch = rob_io_branch_info_bits_is_branch; // @[Exu.scala 46:22]
  assign io_ex_branch_info_o_bits_is_taken = rob_io_branch_info_bits_is_taken; // @[Exu.scala 46:22]
  assign io_ex_branch_info_o_bits_predict_miss = rob_io_branch_info_bits_predict_miss; // @[Exu.scala 46:22]
  assign io_dcache_io_read_req_valid = dcache_io_io_read_req_valid; // @[Exu.scala 51:25]
  assign io_dcache_io_read_req_bits_addr = dcache_io_io_read_req_bits_addr; // @[Exu.scala 51:25]
  assign io_dcache_io_read_req_bits_rob_idx = dcache_io_io_read_req_bits_rob_idx; // @[Exu.scala 51:25]
  assign io_dcache_io_write_req_valid = dcache_io_io_write_req_valid; // @[Exu.scala 53:25]
  assign io_dcache_io_write_req_bits_addr = dcache_io_io_write_req_bits_addr; // @[Exu.scala 53:25]
  assign io_dcache_io_write_req_bits_data = dcache_io_io_write_req_bits_data; // @[Exu.scala 53:25]
  assign io_dcache_io_write_req_bits_byte_mask = dcache_io_io_write_req_bits_byte_mask; // @[Exu.scala 53:25]
  assign io_need_flush = rob_io_need_flush; // @[Exu.scala 55:20]
  assign io_rob_commit_0_valid = rob_io_rob_commit_0_valid; // @[Exu.scala 84:20]
  assign io_rob_commit_0_bits_des_rob = rob_io_rob_commit_0_bits_des_rob; // @[Exu.scala 84:20]
  assign io_rob_commit_1_valid = rob_io_rob_commit_1_valid; // @[Exu.scala 84:20]
  assign io_rob_commit_1_bits_des_rob = rob_io_rob_commit_1_bits_des_rob; // @[Exu.scala 84:20]
  assign decode_clock = clock;
  assign decode_reset = reset;
  assign decode_io_fb_inst_bank_valid = io_fb_inst_bank_i_valid; // @[Exu.scala 37:20]
  assign decode_io_fb_inst_bank_bits_data_0_inst = io_fb_inst_bank_i_bits_data_0_inst; // @[Exu.scala 37:20]
  assign decode_io_fb_inst_bank_bits_data_0_inst_addr = io_fb_inst_bank_i_bits_data_0_inst_addr; // @[Exu.scala 37:20]
  assign decode_io_fb_inst_bank_bits_data_0_gh_backup = io_fb_inst_bank_i_bits_data_0_gh_backup; // @[Exu.scala 37:20]
  assign decode_io_fb_inst_bank_bits_data_0_is_valid = io_fb_inst_bank_i_bits_data_0_is_valid; // @[Exu.scala 37:20]
  assign decode_io_fb_inst_bank_bits_data_0_predict_taken = io_fb_inst_bank_i_bits_data_0_predict_taken; // @[Exu.scala 37:20]
  assign decode_io_fb_inst_bank_bits_data_1_inst = io_fb_inst_bank_i_bits_data_1_inst; // @[Exu.scala 37:20]
  assign decode_io_fb_inst_bank_bits_data_1_inst_addr = io_fb_inst_bank_i_bits_data_1_inst_addr; // @[Exu.scala 37:20]
  assign decode_io_fb_inst_bank_bits_data_1_gh_backup = io_fb_inst_bank_i_bits_data_1_gh_backup; // @[Exu.scala 37:20]
  assign decode_io_fb_inst_bank_bits_data_1_is_valid = io_fb_inst_bank_i_bits_data_1_is_valid; // @[Exu.scala 37:20]
  assign decode_io_fb_inst_bank_bits_data_1_predict_taken = io_fb_inst_bank_i_bits_data_1_predict_taken; // @[Exu.scala 37:20]
  assign decode_io_rob_allocate_allocate_resp_valid = rob_io_rob_allocate_allocate_resp_valid; // @[Exu.scala 39:22]
  assign decode_io_rob_allocate_allocate_resp_bits_rob_idx_0 = rob_io_rob_allocate_allocate_resp_bits_rob_idx_0; // @[Exu.scala 39:22]
  assign decode_io_rob_allocate_allocate_resp_bits_rob_idx_1 = rob_io_rob_allocate_allocate_resp_bits_rob_idx_1; // @[Exu.scala 39:22]
  assign decode_io_rob_allocate_allocate_resp_bits_enq_valid_mask_0 =
    rob_io_rob_allocate_allocate_resp_bits_enq_valid_mask_0; // @[Exu.scala 39:22]
  assign decode_io_rob_allocate_allocate_resp_bits_enq_valid_mask_1 =
    rob_io_rob_allocate_allocate_resp_bits_enq_valid_mask_1; // @[Exu.scala 39:22]
  assign decode_io_need_flush = rob_io_need_flush; // @[Exu.scala 56:20]
  assign rename_clock = clock;
  assign rename_reset = reset;
  assign rename_io_rename_info_valid = decode_io_rename_info_valid; // @[Exu.scala 40:24]
  assign rename_io_rename_info_bits_0_is_valid = decode_io_rename_info_bits_0_is_valid; // @[Exu.scala 40:24]
  assign rename_io_rename_info_bits_0_op1_addr = decode_io_rename_info_bits_0_op1_addr; // @[Exu.scala 40:24]
  assign rename_io_rename_info_bits_0_op2_addr = decode_io_rename_info_bits_0_op2_addr; // @[Exu.scala 40:24]
  assign rename_io_rename_info_bits_0_des_addr = decode_io_rename_info_bits_0_des_addr; // @[Exu.scala 40:24]
  assign rename_io_rename_info_bits_0_des_rob = decode_io_rename_info_bits_0_des_rob; // @[Exu.scala 40:24]
  assign rename_io_rename_info_bits_1_is_valid = decode_io_rename_info_bits_1_is_valid; // @[Exu.scala 40:24]
  assign rename_io_rename_info_bits_1_op1_addr = decode_io_rename_info_bits_1_op1_addr; // @[Exu.scala 40:24]
  assign rename_io_rename_info_bits_1_op2_addr = decode_io_rename_info_bits_1_op2_addr; // @[Exu.scala 40:24]
  assign rename_io_rename_info_bits_1_des_addr = decode_io_rename_info_bits_1_des_addr; // @[Exu.scala 40:24]
  assign rename_io_rename_info_bits_1_des_rob = decode_io_rename_info_bits_1_des_rob; // @[Exu.scala 40:24]
  assign rename_io_rob_commit_0_valid = rob_io_rob_commit_0_valid; // @[Exu.scala 43:23]
  assign rename_io_rob_commit_0_bits_des_rob = rob_io_rob_commit_0_bits_des_rob; // @[Exu.scala 43:23]
  assign rename_io_rob_commit_0_bits_commit_addr = rob_io_rob_commit_0_bits_commit_addr; // @[Exu.scala 43:23]
  assign rename_io_rob_commit_1_valid = rob_io_rob_commit_1_valid; // @[Exu.scala 43:23]
  assign rename_io_rob_commit_1_bits_des_rob = rob_io_rob_commit_1_bits_des_rob; // @[Exu.scala 43:23]
  assign rename_io_rob_commit_1_bits_commit_addr = rob_io_rob_commit_1_bits_commit_addr; // @[Exu.scala 43:23]
  assign rename_io_reg_read_0_op1_data = regfile_io_reg_read_0_op1_data; // @[Exu.scala 41:21]
  assign rename_io_reg_read_0_op2_data = regfile_io_reg_read_0_op2_data; // @[Exu.scala 41:21]
  assign rename_io_reg_read_1_op1_data = regfile_io_reg_read_1_op1_data; // @[Exu.scala 41:21]
  assign rename_io_reg_read_1_op2_data = regfile_io_reg_read_1_op2_data; // @[Exu.scala 41:21]
  assign rename_io_need_flush = rob_io_need_flush; // @[Exu.scala 57:20]
  assign regfile_clock = clock;
  assign regfile_reset = reset;
  assign regfile_io_reg_read_0_op1_addr = rename_io_reg_read_0_op1_addr; // @[Exu.scala 41:21]
  assign regfile_io_reg_read_0_op2_addr = rename_io_reg_read_0_op2_addr; // @[Exu.scala 41:21]
  assign regfile_io_reg_read_1_op1_addr = rename_io_reg_read_1_op1_addr; // @[Exu.scala 41:21]
  assign regfile_io_reg_read_1_op2_addr = rename_io_reg_read_1_op2_addr; // @[Exu.scala 41:21]
  assign regfile_io_rob_commit_i_0_valid = rob_io_rob_commit_0_valid; // @[Exu.scala 45:26]
  assign regfile_io_rob_commit_i_0_bits_commit_addr = rob_io_rob_commit_0_bits_commit_addr; // @[Exu.scala 45:26]
  assign regfile_io_rob_commit_i_0_bits_commit_data = rob_io_rob_commit_0_bits_commit_data; // @[Exu.scala 45:26]
  assign regfile_io_rob_commit_i_1_valid = rob_io_rob_commit_1_valid; // @[Exu.scala 45:26]
  assign regfile_io_rob_commit_i_1_bits_commit_addr = rob_io_rob_commit_1_bits_commit_addr; // @[Exu.scala 45:26]
  assign regfile_io_rob_commit_i_1_bits_commit_data = rob_io_rob_commit_1_bits_commit_data; // @[Exu.scala 45:26]
  assign rob_clock = clock;
  assign rob_reset = reset;
  assign rob_io_rob_allocate_allocate_req_valid = decode_io_rob_allocate_allocate_req_valid; // @[Exu.scala 39:22]
  assign rob_io_rob_allocate_allocate_req_bits_0 = decode_io_rob_allocate_allocate_req_bits_0; // @[Exu.scala 39:22]
  assign rob_io_rob_allocate_allocate_req_bits_1 = decode_io_rob_allocate_allocate_req_bits_1; // @[Exu.scala 39:22]
  assign rob_io_rob_allocate_allocate_info_valid = decode_io_rob_allocate_allocate_info_valid; // @[Exu.scala 39:22]
  assign rob_io_rob_allocate_allocate_info_bits_0_rob_idx = decode_io_rob_allocate_allocate_info_bits_0_rob_idx; // @[Exu.scala 39:22]
  assign rob_io_rob_allocate_allocate_info_bits_0_inst_valid = decode_io_rob_allocate_allocate_info_bits_0_inst_valid; // @[Exu.scala 39:22]
  assign rob_io_rob_allocate_allocate_info_bits_0_inst_addr = decode_io_rob_allocate_allocate_info_bits_0_inst_addr; // @[Exu.scala 39:22]
  assign rob_io_rob_allocate_allocate_info_bits_0_uop = decode_io_rob_allocate_allocate_info_bits_0_uop; // @[Exu.scala 39:22]
  assign rob_io_rob_allocate_allocate_info_bits_0_unit_sel = decode_io_rob_allocate_allocate_info_bits_0_unit_sel; // @[Exu.scala 39:22]
  assign rob_io_rob_allocate_allocate_info_bits_0_need_imm = decode_io_rob_allocate_allocate_info_bits_0_need_imm; // @[Exu.scala 39:22]
  assign rob_io_rob_allocate_allocate_info_bits_0_commit_addr = decode_io_rob_allocate_allocate_info_bits_0_commit_addr; // @[Exu.scala 39:22]
  assign rob_io_rob_allocate_allocate_info_bits_0_gh_info = decode_io_rob_allocate_allocate_info_bits_0_gh_info; // @[Exu.scala 39:22]
  assign rob_io_rob_allocate_allocate_info_bits_0_imm_data = decode_io_rob_allocate_allocate_info_bits_0_imm_data; // @[Exu.scala 39:22]
  assign rob_io_rob_allocate_allocate_info_bits_0_flush_on_commit =
    decode_io_rob_allocate_allocate_info_bits_0_flush_on_commit; // @[Exu.scala 39:22]
  assign rob_io_rob_allocate_allocate_info_bits_0_predict_taken =
    decode_io_rob_allocate_allocate_info_bits_0_predict_taken; // @[Exu.scala 39:22]
  assign rob_io_rob_allocate_allocate_info_bits_1_rob_idx = decode_io_rob_allocate_allocate_info_bits_1_rob_idx; // @[Exu.scala 39:22]
  assign rob_io_rob_allocate_allocate_info_bits_1_inst_valid = decode_io_rob_allocate_allocate_info_bits_1_inst_valid; // @[Exu.scala 39:22]
  assign rob_io_rob_allocate_allocate_info_bits_1_inst_addr = decode_io_rob_allocate_allocate_info_bits_1_inst_addr; // @[Exu.scala 39:22]
  assign rob_io_rob_allocate_allocate_info_bits_1_uop = decode_io_rob_allocate_allocate_info_bits_1_uop; // @[Exu.scala 39:22]
  assign rob_io_rob_allocate_allocate_info_bits_1_unit_sel = decode_io_rob_allocate_allocate_info_bits_1_unit_sel; // @[Exu.scala 39:22]
  assign rob_io_rob_allocate_allocate_info_bits_1_need_imm = decode_io_rob_allocate_allocate_info_bits_1_need_imm; // @[Exu.scala 39:22]
  assign rob_io_rob_allocate_allocate_info_bits_1_commit_addr = decode_io_rob_allocate_allocate_info_bits_1_commit_addr; // @[Exu.scala 39:22]
  assign rob_io_rob_allocate_allocate_info_bits_1_gh_info = decode_io_rob_allocate_allocate_info_bits_1_gh_info; // @[Exu.scala 39:22]
  assign rob_io_rob_allocate_allocate_info_bits_1_imm_data = decode_io_rob_allocate_allocate_info_bits_1_imm_data; // @[Exu.scala 39:22]
  assign rob_io_rob_allocate_allocate_info_bits_1_flush_on_commit =
    decode_io_rob_allocate_allocate_info_bits_1_flush_on_commit; // @[Exu.scala 39:22]
  assign rob_io_rob_allocate_allocate_info_bits_1_predict_taken =
    decode_io_rob_allocate_allocate_info_bits_1_predict_taken; // @[Exu.scala 39:22]
  assign rob_io_rob_init_info_valid = rename_io_rob_init_info_valid; // @[Exu.scala 42:23]
  assign rob_io_rob_init_info_bits_0_is_valid = rename_io_rob_init_info_bits_0_is_valid; // @[Exu.scala 42:23]
  assign rob_io_rob_init_info_bits_0_des_rob = rename_io_rob_init_info_bits_0_des_rob; // @[Exu.scala 42:23]
  assign rob_io_rob_init_info_bits_0_op1_rob = rename_io_rob_init_info_bits_0_op1_rob; // @[Exu.scala 42:23]
  assign rob_io_rob_init_info_bits_0_op2_rob = rename_io_rob_init_info_bits_0_op2_rob; // @[Exu.scala 42:23]
  assign rob_io_rob_init_info_bits_0_op1_regData = rename_io_rob_init_info_bits_0_op1_regData; // @[Exu.scala 42:23]
  assign rob_io_rob_init_info_bits_0_op2_regData = rename_io_rob_init_info_bits_0_op2_regData; // @[Exu.scala 42:23]
  assign rob_io_rob_init_info_bits_0_op1_in_rob = rename_io_rob_init_info_bits_0_op1_in_rob; // @[Exu.scala 42:23]
  assign rob_io_rob_init_info_bits_0_op2_in_rob = rename_io_rob_init_info_bits_0_op2_in_rob; // @[Exu.scala 42:23]
  assign rob_io_rob_init_info_bits_1_is_valid = rename_io_rob_init_info_bits_1_is_valid; // @[Exu.scala 42:23]
  assign rob_io_rob_init_info_bits_1_des_rob = rename_io_rob_init_info_bits_1_des_rob; // @[Exu.scala 42:23]
  assign rob_io_rob_init_info_bits_1_op1_rob = rename_io_rob_init_info_bits_1_op1_rob; // @[Exu.scala 42:23]
  assign rob_io_rob_init_info_bits_1_op2_rob = rename_io_rob_init_info_bits_1_op2_rob; // @[Exu.scala 42:23]
  assign rob_io_rob_init_info_bits_1_op1_regData = rename_io_rob_init_info_bits_1_op1_regData; // @[Exu.scala 42:23]
  assign rob_io_rob_init_info_bits_1_op2_regData = rename_io_rob_init_info_bits_1_op2_regData; // @[Exu.scala 42:23]
  assign rob_io_rob_init_info_bits_1_op1_in_rob = rename_io_rob_init_info_bits_1_op1_in_rob; // @[Exu.scala 42:23]
  assign rob_io_rob_init_info_bits_1_op2_in_rob = rename_io_rob_init_info_bits_1_op2_in_rob; // @[Exu.scala 42:23]
  assign rob_io_wb_info_i_0_valid = alu0_io_wb_info_valid; // @[Exu.scala 67:22]
  assign rob_io_wb_info_i_0_bits_rob_idx = alu0_io_wb_info_bits_rob_idx; // @[Exu.scala 67:22]
  assign rob_io_wb_info_i_0_bits_data = alu0_io_wb_info_bits_data; // @[Exu.scala 67:22]
  assign rob_io_wb_info_i_1_valid = alu1_io_wb_info_valid; // @[Exu.scala 68:22]
  assign rob_io_wb_info_i_1_bits_rob_idx = alu1_io_wb_info_bits_rob_idx; // @[Exu.scala 68:22]
  assign rob_io_wb_info_i_1_bits_data = alu1_io_wb_info_bits_data; // @[Exu.scala 68:22]
  assign rob_io_wb_info_i_2_valid = bju0_io_wb_info_valid; // @[Exu.scala 70:22]
  assign rob_io_wb_info_i_2_bits_rob_idx = bju0_io_wb_info_bits_rob_idx; // @[Exu.scala 70:22]
  assign rob_io_wb_info_i_2_bits_data = bju0_io_wb_info_bits_data; // @[Exu.scala 70:22]
  assign rob_io_wb_info_i_2_bits_target_addr = bju0_io_wb_info_bits_target_addr; // @[Exu.scala 70:22]
  assign rob_io_wb_info_i_2_bits_is_taken = bju0_io_wb_info_bits_is_taken; // @[Exu.scala 70:22]
  assign rob_io_wb_info_i_2_bits_predict_miss = bju0_io_wb_info_bits_predict_miss; // @[Exu.scala 70:22]
  assign rob_io_wb_info_i_3_valid = mdu_io_wb_info_valid; // @[Exu.scala 72:22]
  assign rob_io_wb_info_i_3_bits_rob_idx = mdu_io_wb_info_bits_rob_idx; // @[Exu.scala 72:22]
  assign rob_io_wb_info_i_3_bits_data = mdu_io_wb_info_bits_data; // @[Exu.scala 72:22]
  assign rob_io_wb_info_i_4_valid = lsu_io_wb_info_valid; // @[Exu.scala 73:22]
  assign rob_io_wb_info_i_4_bits_rob_idx = lsu_io_wb_info_bits_rob_idx; // @[Exu.scala 73:22]
  assign rob_io_wb_info_i_4_bits_data = lsu_io_wb_info_bits_data; // @[Exu.scala 73:22]
  assign rob_io_dispatch_info_o_4_ready = lsu_io_dispatch_info_ready; // @[Exu.scala 81:28]
  assign alu0_clock = clock;
  assign alu0_reset = reset;
  assign alu0_io_dispatch_info_valid = rob_io_dispatch_info_o_0_valid; // @[Exu.scala 75:28]
  assign alu0_io_dispatch_info_bits_uop = rob_io_dispatch_info_o_0_bits_uop; // @[Exu.scala 75:28]
  assign alu0_io_dispatch_info_bits_need_imm = rob_io_dispatch_info_o_0_bits_need_imm; // @[Exu.scala 75:28]
  assign alu0_io_dispatch_info_bits_rob_idx = rob_io_dispatch_info_o_0_bits_rob_idx; // @[Exu.scala 75:28]
  assign alu0_io_dispatch_info_bits_op1_data = rob_io_dispatch_info_o_0_bits_op1_data; // @[Exu.scala 75:28]
  assign alu0_io_dispatch_info_bits_op2_data = rob_io_dispatch_info_o_0_bits_op2_data; // @[Exu.scala 75:28]
  assign alu0_io_dispatch_info_bits_imm_data = rob_io_dispatch_info_o_0_bits_imm_data; // @[Exu.scala 75:28]
  assign alu0_io_need_flush = rob_io_need_flush; // @[Exu.scala 58:20]
  assign alu1_clock = clock;
  assign alu1_reset = reset;
  assign alu1_io_dispatch_info_valid = rob_io_dispatch_info_o_1_valid; // @[Exu.scala 76:28]
  assign alu1_io_dispatch_info_bits_uop = rob_io_dispatch_info_o_1_bits_uop; // @[Exu.scala 76:28]
  assign alu1_io_dispatch_info_bits_need_imm = rob_io_dispatch_info_o_1_bits_need_imm; // @[Exu.scala 76:28]
  assign alu1_io_dispatch_info_bits_rob_idx = rob_io_dispatch_info_o_1_bits_rob_idx; // @[Exu.scala 76:28]
  assign alu1_io_dispatch_info_bits_op1_data = rob_io_dispatch_info_o_1_bits_op1_data; // @[Exu.scala 76:28]
  assign alu1_io_dispatch_info_bits_op2_data = rob_io_dispatch_info_o_1_bits_op2_data; // @[Exu.scala 76:28]
  assign alu1_io_dispatch_info_bits_imm_data = rob_io_dispatch_info_o_1_bits_imm_data; // @[Exu.scala 76:28]
  assign alu1_io_need_flush = rob_io_need_flush; // @[Exu.scala 59:20]
  assign bju0_clock = clock;
  assign bju0_reset = reset;
  assign bju0_io_dispatch_info_valid = rob_io_dispatch_info_o_2_valid; // @[Exu.scala 78:28]
  assign bju0_io_dispatch_info_bits_uop = rob_io_dispatch_info_o_2_bits_uop; // @[Exu.scala 78:28]
  assign bju0_io_dispatch_info_bits_rob_idx = rob_io_dispatch_info_o_2_bits_rob_idx; // @[Exu.scala 78:28]
  assign bju0_io_dispatch_info_bits_inst_addr = rob_io_dispatch_info_o_2_bits_inst_addr; // @[Exu.scala 78:28]
  assign bju0_io_dispatch_info_bits_op1_data = rob_io_dispatch_info_o_2_bits_op1_data; // @[Exu.scala 78:28]
  assign bju0_io_dispatch_info_bits_op2_data = rob_io_dispatch_info_o_2_bits_op2_data; // @[Exu.scala 78:28]
  assign bju0_io_dispatch_info_bits_imm_data = rob_io_dispatch_info_o_2_bits_imm_data; // @[Exu.scala 78:28]
  assign bju0_io_dispatch_info_bits_predict_taken = rob_io_dispatch_info_o_2_bits_predict_taken; // @[Exu.scala 78:28]
  assign bju0_io_need_flush = rob_io_need_flush; // @[Exu.scala 61:20]
  assign lsu_clock = clock;
  assign lsu_reset = reset;
  assign lsu_io_dispatch_info_valid = rob_io_dispatch_info_o_4_valid; // @[Exu.scala 81:28]
  assign lsu_io_dispatch_info_bits_uop = rob_io_dispatch_info_o_4_bits_uop; // @[Exu.scala 81:28]
  assign lsu_io_dispatch_info_bits_rob_idx = rob_io_dispatch_info_o_4_bits_rob_idx; // @[Exu.scala 81:28]
  assign lsu_io_dispatch_info_bits_op1_data = rob_io_dispatch_info_o_4_bits_op1_data; // @[Exu.scala 81:28]
  assign lsu_io_dispatch_info_bits_op2_data = rob_io_dispatch_info_o_4_bits_op2_data; // @[Exu.scala 81:28]
  assign lsu_io_dispatch_info_bits_imm_data = rob_io_dispatch_info_o_4_bits_imm_data; // @[Exu.scala 81:28]
  assign lsu_io_rob_commit_0_valid = rob_io_rob_commit_0_valid; // @[Exu.scala 47:20]
  assign lsu_io_rob_commit_0_bits_des_rob = rob_io_rob_commit_0_bits_des_rob; // @[Exu.scala 47:20]
  assign lsu_io_rob_commit_1_valid = rob_io_rob_commit_1_valid; // @[Exu.scala 47:20]
  assign lsu_io_rob_commit_1_bits_des_rob = rob_io_rob_commit_1_bits_des_rob; // @[Exu.scala 47:20]
  assign lsu_io_cache_read_ready = dcache_io_dcache_read_req_ready; // @[Exu.scala 48:21]
  assign lsu_io_cache_write_ready = dcache_io_dcache_write_req_ready; // @[Exu.scala 49:21]
  assign lsu_io_cache_resp_data = dcache_io_dcache_read_resp_data; // @[Exu.scala 50:21]
  assign lsu_io_need_flush = rob_io_need_flush; // @[Exu.scala 63:20]
  assign mdu_clock = clock;
  assign mdu_reset = reset;
  assign mdu_io_dispatch_info_valid = rob_io_dispatch_info_o_3_valid; // @[Exu.scala 80:28]
  assign mdu_io_dispatch_info_bits_rob_idx = rob_io_dispatch_info_o_3_bits_rob_idx; // @[Exu.scala 80:28]
  assign mdu_io_dispatch_info_bits_op1_data = rob_io_dispatch_info_o_3_bits_op1_data; // @[Exu.scala 80:28]
  assign mdu_io_dispatch_info_bits_op2_data = rob_io_dispatch_info_o_3_bits_op2_data; // @[Exu.scala 80:28]
  assign mdu_io_need_flush = rob_io_need_flush; // @[Exu.scala 64:20]
  assign dcache_io_dcache_read_req_valid = lsu_io_cache_read_valid; // @[Exu.scala 48:21]
  assign dcache_io_dcache_read_req_bits_addr = lsu_io_cache_read_bits_addr; // @[Exu.scala 48:21]
  assign dcache_io_dcache_read_req_bits_rob_idx = lsu_io_cache_read_bits_rob_idx; // @[Exu.scala 48:21]
  assign dcache_io_dcache_write_req_valid = lsu_io_cache_write_valid; // @[Exu.scala 49:21]
  assign dcache_io_dcache_write_req_bits_addr = lsu_io_cache_write_bits_addr; // @[Exu.scala 49:21]
  assign dcache_io_dcache_write_req_bits_data = lsu_io_cache_write_bits_data; // @[Exu.scala 49:21]
  assign dcache_io_dcache_write_req_bits_byte_mask = lsu_io_cache_write_bits_byte_mask; // @[Exu.scala 49:21]
  assign dcache_io_io_read_req_ready = io_dcache_io_read_req_ready; // @[Exu.scala 51:25]
  assign dcache_io_io_read_resp_bits_data = io_dcache_io_read_resp_bits_data; // @[Exu.scala 52:25]
  assign dcache_io_io_write_req_ready = io_dcache_io_write_req_ready; // @[Exu.scala 53:25]
endmodule
module Core(
  input          clock,
  input          reset,
  input          io_icache_io_read_req_ready,
  output         io_icache_io_read_req_valid,
  output [31:0]  io_icache_io_read_req_bits_addr,
  input  [255:0] io_icache_io_read_resp_bits_data,
  input          io_dcache_io_read_req_ready,
  output         io_dcache_io_read_req_valid,
  output [31:0]  io_dcache_io_read_req_bits_addr,
  output [3:0]   io_dcache_io_read_req_bits_rob_idx,
  input  [31:0]  io_dcache_io_read_resp_bits_data,
  input          io_dcache_io_write_req_ready,
  output         io_dcache_io_write_req_valid,
  output [31:0]  io_dcache_io_write_req_bits_addr,
  output [31:0]  io_dcache_io_write_req_bits_data,
  output [3:0]   io_dcache_io_write_req_bits_byte_mask,
  output         io_need_flush,
  output         io_rob_commit_0_valid,
  output [2:0]   io_rob_commit_0_bits_des_rob,
  output         io_rob_commit_1_valid,
  output [2:0]   io_rob_commit_1_bits_des_rob,
  output         io_icache_debug_state,
  output         io_icache_debug_hit_cache,
  output         io_icache_debug_cache_we,
  output [19:0]  io_icache_debug_cache_read_tag,
  output         io_icache_debug_icache_req_valid,
  output [31:0]  io_icache_debug_icache_req_bits_addr,
  output [7:0]   io_bpu_debug_branch_mask,
  output [7:0]   io_bpu_debug_fetched_mask,
  output [7:0]   io_bpu_debug_predict_branch,
  output [31:0]  io_bpu_debug_predict_addr,
  output         io_bpu_debug_is_taken,
  output         io_bpu_debug_take_delay,
  output [31:0]  io_bpu_debug_inst_packet_0,
  output [31:0]  io_bpu_debug_inst_packet_1,
  output [31:0]  io_bpu_debug_inst_packet_2,
  output [31:0]  io_bpu_debug_inst_packet_3,
  output [31:0]  io_bpu_debug_inst_packet_4,
  output [31:0]  io_bpu_debug_inst_packet_5,
  output [31:0]  io_bpu_debug_inst_packet_6,
  output [31:0]  io_bpu_debug_inst_packet_7
);
  wire  ifu_clock; // @[Core.scala 25:19]
  wire  ifu_reset; // @[Core.scala 25:19]
  wire  ifu_io_ex_branch_info_i_valid; // @[Core.scala 25:19]
  wire [31:0] ifu_io_ex_branch_info_i_bits_target_addr; // @[Core.scala 25:19]
  wire [31:0] ifu_io_ex_branch_info_i_bits_inst_addr; // @[Core.scala 25:19]
  wire [3:0] ifu_io_ex_branch_info_i_bits_gh_update; // @[Core.scala 25:19]
  wire  ifu_io_ex_branch_info_i_bits_is_branch; // @[Core.scala 25:19]
  wire  ifu_io_ex_branch_info_i_bits_is_taken; // @[Core.scala 25:19]
  wire  ifu_io_ex_branch_info_i_bits_predict_miss; // @[Core.scala 25:19]
  wire  ifu_io_fb_inst_bank_o_valid; // @[Core.scala 25:19]
  wire [31:0] ifu_io_fb_inst_bank_o_bits_data_0_inst; // @[Core.scala 25:19]
  wire [31:0] ifu_io_fb_inst_bank_o_bits_data_0_inst_addr; // @[Core.scala 25:19]
  wire [3:0] ifu_io_fb_inst_bank_o_bits_data_0_gh_backup; // @[Core.scala 25:19]
  wire  ifu_io_fb_inst_bank_o_bits_data_0_is_valid; // @[Core.scala 25:19]
  wire  ifu_io_fb_inst_bank_o_bits_data_0_predict_taken; // @[Core.scala 25:19]
  wire [31:0] ifu_io_fb_inst_bank_o_bits_data_1_inst; // @[Core.scala 25:19]
  wire [31:0] ifu_io_fb_inst_bank_o_bits_data_1_inst_addr; // @[Core.scala 25:19]
  wire [3:0] ifu_io_fb_inst_bank_o_bits_data_1_gh_backup; // @[Core.scala 25:19]
  wire  ifu_io_fb_inst_bank_o_bits_data_1_is_valid; // @[Core.scala 25:19]
  wire  ifu_io_fb_inst_bank_o_bits_data_1_predict_taken; // @[Core.scala 25:19]
  wire  ifu_io_fb_resp_deq_valid_0; // @[Core.scala 25:19]
  wire  ifu_io_fb_resp_deq_valid_1; // @[Core.scala 25:19]
  wire  ifu_io_icache_io_read_req_ready; // @[Core.scala 25:19]
  wire  ifu_io_icache_io_read_req_valid; // @[Core.scala 25:19]
  wire [31:0] ifu_io_icache_io_read_req_bits_addr; // @[Core.scala 25:19]
  wire [255:0] ifu_io_icache_io_read_resp_bits_data; // @[Core.scala 25:19]
  wire  ifu_io_icache_debug_state; // @[Core.scala 25:19]
  wire  ifu_io_icache_debug_hit_cache; // @[Core.scala 25:19]
  wire  ifu_io_icache_debug_cache_we; // @[Core.scala 25:19]
  wire [19:0] ifu_io_icache_debug_cache_read_tag; // @[Core.scala 25:19]
  wire  ifu_io_icache_debug_icache_req_valid; // @[Core.scala 25:19]
  wire [31:0] ifu_io_icache_debug_icache_req_bits_addr; // @[Core.scala 25:19]
  wire [7:0] ifu_io_bpu_debug_branch_mask; // @[Core.scala 25:19]
  wire [7:0] ifu_io_bpu_debug_fetched_mask; // @[Core.scala 25:19]
  wire [7:0] ifu_io_bpu_debug_predict_branch; // @[Core.scala 25:19]
  wire [31:0] ifu_io_bpu_debug_predict_addr; // @[Core.scala 25:19]
  wire  ifu_io_bpu_debug_is_taken; // @[Core.scala 25:19]
  wire  ifu_io_bpu_debug_take_delay; // @[Core.scala 25:19]
  wire [31:0] ifu_io_bpu_debug_inst_packet_0; // @[Core.scala 25:19]
  wire [31:0] ifu_io_bpu_debug_inst_packet_1; // @[Core.scala 25:19]
  wire [31:0] ifu_io_bpu_debug_inst_packet_2; // @[Core.scala 25:19]
  wire [31:0] ifu_io_bpu_debug_inst_packet_3; // @[Core.scala 25:19]
  wire [31:0] ifu_io_bpu_debug_inst_packet_4; // @[Core.scala 25:19]
  wire [31:0] ifu_io_bpu_debug_inst_packet_5; // @[Core.scala 25:19]
  wire [31:0] ifu_io_bpu_debug_inst_packet_6; // @[Core.scala 25:19]
  wire [31:0] ifu_io_bpu_debug_inst_packet_7; // @[Core.scala 25:19]
  wire  exu_clock; // @[Core.scala 26:19]
  wire  exu_reset; // @[Core.scala 26:19]
  wire  exu_io_fb_inst_bank_i_valid; // @[Core.scala 26:19]
  wire [31:0] exu_io_fb_inst_bank_i_bits_data_0_inst; // @[Core.scala 26:19]
  wire [31:0] exu_io_fb_inst_bank_i_bits_data_0_inst_addr; // @[Core.scala 26:19]
  wire [3:0] exu_io_fb_inst_bank_i_bits_data_0_gh_backup; // @[Core.scala 26:19]
  wire  exu_io_fb_inst_bank_i_bits_data_0_is_valid; // @[Core.scala 26:19]
  wire  exu_io_fb_inst_bank_i_bits_data_0_predict_taken; // @[Core.scala 26:19]
  wire [31:0] exu_io_fb_inst_bank_i_bits_data_1_inst; // @[Core.scala 26:19]
  wire [31:0] exu_io_fb_inst_bank_i_bits_data_1_inst_addr; // @[Core.scala 26:19]
  wire [3:0] exu_io_fb_inst_bank_i_bits_data_1_gh_backup; // @[Core.scala 26:19]
  wire  exu_io_fb_inst_bank_i_bits_data_1_is_valid; // @[Core.scala 26:19]
  wire  exu_io_fb_inst_bank_i_bits_data_1_predict_taken; // @[Core.scala 26:19]
  wire  exu_io_fb_resp_deq_valid_0; // @[Core.scala 26:19]
  wire  exu_io_fb_resp_deq_valid_1; // @[Core.scala 26:19]
  wire  exu_io_ex_branch_info_o_valid; // @[Core.scala 26:19]
  wire [31:0] exu_io_ex_branch_info_o_bits_target_addr; // @[Core.scala 26:19]
  wire [31:0] exu_io_ex_branch_info_o_bits_inst_addr; // @[Core.scala 26:19]
  wire [3:0] exu_io_ex_branch_info_o_bits_gh_update; // @[Core.scala 26:19]
  wire  exu_io_ex_branch_info_o_bits_is_branch; // @[Core.scala 26:19]
  wire  exu_io_ex_branch_info_o_bits_is_taken; // @[Core.scala 26:19]
  wire  exu_io_ex_branch_info_o_bits_predict_miss; // @[Core.scala 26:19]
  wire  exu_io_dcache_io_read_req_ready; // @[Core.scala 26:19]
  wire  exu_io_dcache_io_read_req_valid; // @[Core.scala 26:19]
  wire [31:0] exu_io_dcache_io_read_req_bits_addr; // @[Core.scala 26:19]
  wire [3:0] exu_io_dcache_io_read_req_bits_rob_idx; // @[Core.scala 26:19]
  wire [31:0] exu_io_dcache_io_read_resp_bits_data; // @[Core.scala 26:19]
  wire  exu_io_dcache_io_write_req_ready; // @[Core.scala 26:19]
  wire  exu_io_dcache_io_write_req_valid; // @[Core.scala 26:19]
  wire [31:0] exu_io_dcache_io_write_req_bits_addr; // @[Core.scala 26:19]
  wire [31:0] exu_io_dcache_io_write_req_bits_data; // @[Core.scala 26:19]
  wire [3:0] exu_io_dcache_io_write_req_bits_byte_mask; // @[Core.scala 26:19]
  wire  exu_io_need_flush; // @[Core.scala 26:19]
  wire  exu_io_rob_commit_0_valid; // @[Core.scala 26:19]
  wire [2:0] exu_io_rob_commit_0_bits_des_rob; // @[Core.scala 26:19]
  wire  exu_io_rob_commit_1_valid; // @[Core.scala 26:19]
  wire [2:0] exu_io_rob_commit_1_bits_des_rob; // @[Core.scala 26:19]
  Ifu ifu ( // @[Core.scala 25:19]
    .clock(ifu_clock),
    .reset(ifu_reset),
    .io_ex_branch_info_i_valid(ifu_io_ex_branch_info_i_valid),
    .io_ex_branch_info_i_bits_target_addr(ifu_io_ex_branch_info_i_bits_target_addr),
    .io_ex_branch_info_i_bits_inst_addr(ifu_io_ex_branch_info_i_bits_inst_addr),
    .io_ex_branch_info_i_bits_gh_update(ifu_io_ex_branch_info_i_bits_gh_update),
    .io_ex_branch_info_i_bits_is_branch(ifu_io_ex_branch_info_i_bits_is_branch),
    .io_ex_branch_info_i_bits_is_taken(ifu_io_ex_branch_info_i_bits_is_taken),
    .io_ex_branch_info_i_bits_predict_miss(ifu_io_ex_branch_info_i_bits_predict_miss),
    .io_fb_inst_bank_o_valid(ifu_io_fb_inst_bank_o_valid),
    .io_fb_inst_bank_o_bits_data_0_inst(ifu_io_fb_inst_bank_o_bits_data_0_inst),
    .io_fb_inst_bank_o_bits_data_0_inst_addr(ifu_io_fb_inst_bank_o_bits_data_0_inst_addr),
    .io_fb_inst_bank_o_bits_data_0_gh_backup(ifu_io_fb_inst_bank_o_bits_data_0_gh_backup),
    .io_fb_inst_bank_o_bits_data_0_is_valid(ifu_io_fb_inst_bank_o_bits_data_0_is_valid),
    .io_fb_inst_bank_o_bits_data_0_predict_taken(ifu_io_fb_inst_bank_o_bits_data_0_predict_taken),
    .io_fb_inst_bank_o_bits_data_1_inst(ifu_io_fb_inst_bank_o_bits_data_1_inst),
    .io_fb_inst_bank_o_bits_data_1_inst_addr(ifu_io_fb_inst_bank_o_bits_data_1_inst_addr),
    .io_fb_inst_bank_o_bits_data_1_gh_backup(ifu_io_fb_inst_bank_o_bits_data_1_gh_backup),
    .io_fb_inst_bank_o_bits_data_1_is_valid(ifu_io_fb_inst_bank_o_bits_data_1_is_valid),
    .io_fb_inst_bank_o_bits_data_1_predict_taken(ifu_io_fb_inst_bank_o_bits_data_1_predict_taken),
    .io_fb_resp_deq_valid_0(ifu_io_fb_resp_deq_valid_0),
    .io_fb_resp_deq_valid_1(ifu_io_fb_resp_deq_valid_1),
    .io_icache_io_read_req_ready(ifu_io_icache_io_read_req_ready),
    .io_icache_io_read_req_valid(ifu_io_icache_io_read_req_valid),
    .io_icache_io_read_req_bits_addr(ifu_io_icache_io_read_req_bits_addr),
    .io_icache_io_read_resp_bits_data(ifu_io_icache_io_read_resp_bits_data),
    .io_icache_debug_state(ifu_io_icache_debug_state),
    .io_icache_debug_hit_cache(ifu_io_icache_debug_hit_cache),
    .io_icache_debug_cache_we(ifu_io_icache_debug_cache_we),
    .io_icache_debug_cache_read_tag(ifu_io_icache_debug_cache_read_tag),
    .io_icache_debug_icache_req_valid(ifu_io_icache_debug_icache_req_valid),
    .io_icache_debug_icache_req_bits_addr(ifu_io_icache_debug_icache_req_bits_addr),
    .io_bpu_debug_branch_mask(ifu_io_bpu_debug_branch_mask),
    .io_bpu_debug_fetched_mask(ifu_io_bpu_debug_fetched_mask),
    .io_bpu_debug_predict_branch(ifu_io_bpu_debug_predict_branch),
    .io_bpu_debug_predict_addr(ifu_io_bpu_debug_predict_addr),
    .io_bpu_debug_is_taken(ifu_io_bpu_debug_is_taken),
    .io_bpu_debug_take_delay(ifu_io_bpu_debug_take_delay),
    .io_bpu_debug_inst_packet_0(ifu_io_bpu_debug_inst_packet_0),
    .io_bpu_debug_inst_packet_1(ifu_io_bpu_debug_inst_packet_1),
    .io_bpu_debug_inst_packet_2(ifu_io_bpu_debug_inst_packet_2),
    .io_bpu_debug_inst_packet_3(ifu_io_bpu_debug_inst_packet_3),
    .io_bpu_debug_inst_packet_4(ifu_io_bpu_debug_inst_packet_4),
    .io_bpu_debug_inst_packet_5(ifu_io_bpu_debug_inst_packet_5),
    .io_bpu_debug_inst_packet_6(ifu_io_bpu_debug_inst_packet_6),
    .io_bpu_debug_inst_packet_7(ifu_io_bpu_debug_inst_packet_7)
  );
  Exu exu ( // @[Core.scala 26:19]
    .clock(exu_clock),
    .reset(exu_reset),
    .io_fb_inst_bank_i_valid(exu_io_fb_inst_bank_i_valid),
    .io_fb_inst_bank_i_bits_data_0_inst(exu_io_fb_inst_bank_i_bits_data_0_inst),
    .io_fb_inst_bank_i_bits_data_0_inst_addr(exu_io_fb_inst_bank_i_bits_data_0_inst_addr),
    .io_fb_inst_bank_i_bits_data_0_gh_backup(exu_io_fb_inst_bank_i_bits_data_0_gh_backup),
    .io_fb_inst_bank_i_bits_data_0_is_valid(exu_io_fb_inst_bank_i_bits_data_0_is_valid),
    .io_fb_inst_bank_i_bits_data_0_predict_taken(exu_io_fb_inst_bank_i_bits_data_0_predict_taken),
    .io_fb_inst_bank_i_bits_data_1_inst(exu_io_fb_inst_bank_i_bits_data_1_inst),
    .io_fb_inst_bank_i_bits_data_1_inst_addr(exu_io_fb_inst_bank_i_bits_data_1_inst_addr),
    .io_fb_inst_bank_i_bits_data_1_gh_backup(exu_io_fb_inst_bank_i_bits_data_1_gh_backup),
    .io_fb_inst_bank_i_bits_data_1_is_valid(exu_io_fb_inst_bank_i_bits_data_1_is_valid),
    .io_fb_inst_bank_i_bits_data_1_predict_taken(exu_io_fb_inst_bank_i_bits_data_1_predict_taken),
    .io_fb_resp_deq_valid_0(exu_io_fb_resp_deq_valid_0),
    .io_fb_resp_deq_valid_1(exu_io_fb_resp_deq_valid_1),
    .io_ex_branch_info_o_valid(exu_io_ex_branch_info_o_valid),
    .io_ex_branch_info_o_bits_target_addr(exu_io_ex_branch_info_o_bits_target_addr),
    .io_ex_branch_info_o_bits_inst_addr(exu_io_ex_branch_info_o_bits_inst_addr),
    .io_ex_branch_info_o_bits_gh_update(exu_io_ex_branch_info_o_bits_gh_update),
    .io_ex_branch_info_o_bits_is_branch(exu_io_ex_branch_info_o_bits_is_branch),
    .io_ex_branch_info_o_bits_is_taken(exu_io_ex_branch_info_o_bits_is_taken),
    .io_ex_branch_info_o_bits_predict_miss(exu_io_ex_branch_info_o_bits_predict_miss),
    .io_dcache_io_read_req_ready(exu_io_dcache_io_read_req_ready),
    .io_dcache_io_read_req_valid(exu_io_dcache_io_read_req_valid),
    .io_dcache_io_read_req_bits_addr(exu_io_dcache_io_read_req_bits_addr),
    .io_dcache_io_read_req_bits_rob_idx(exu_io_dcache_io_read_req_bits_rob_idx),
    .io_dcache_io_read_resp_bits_data(exu_io_dcache_io_read_resp_bits_data),
    .io_dcache_io_write_req_ready(exu_io_dcache_io_write_req_ready),
    .io_dcache_io_write_req_valid(exu_io_dcache_io_write_req_valid),
    .io_dcache_io_write_req_bits_addr(exu_io_dcache_io_write_req_bits_addr),
    .io_dcache_io_write_req_bits_data(exu_io_dcache_io_write_req_bits_data),
    .io_dcache_io_write_req_bits_byte_mask(exu_io_dcache_io_write_req_bits_byte_mask),
    .io_need_flush(exu_io_need_flush),
    .io_rob_commit_0_valid(exu_io_rob_commit_0_valid),
    .io_rob_commit_0_bits_des_rob(exu_io_rob_commit_0_bits_des_rob),
    .io_rob_commit_1_valid(exu_io_rob_commit_1_valid),
    .io_rob_commit_1_bits_des_rob(exu_io_rob_commit_1_bits_des_rob)
  );
  assign io_icache_io_read_req_valid = ifu_io_icache_io_read_req_valid; // @[Core.scala 31:24]
  assign io_icache_io_read_req_bits_addr = ifu_io_icache_io_read_req_bits_addr; // @[Core.scala 31:24]
  assign io_dcache_io_read_req_valid = exu_io_dcache_io_read_req_valid; // @[Core.scala 34:25]
  assign io_dcache_io_read_req_bits_addr = exu_io_dcache_io_read_req_bits_addr; // @[Core.scala 34:25]
  assign io_dcache_io_read_req_bits_rob_idx = exu_io_dcache_io_read_req_bits_rob_idx; // @[Core.scala 34:25]
  assign io_dcache_io_write_req_valid = exu_io_dcache_io_write_req_valid; // @[Core.scala 36:25]
  assign io_dcache_io_write_req_bits_addr = exu_io_dcache_io_write_req_bits_addr; // @[Core.scala 36:25]
  assign io_dcache_io_write_req_bits_data = exu_io_dcache_io_write_req_bits_data; // @[Core.scala 36:25]
  assign io_dcache_io_write_req_bits_byte_mask = exu_io_dcache_io_write_req_bits_byte_mask; // @[Core.scala 36:25]
  assign io_need_flush = exu_io_need_flush; // @[Core.scala 38:16]
  assign io_rob_commit_0_valid = exu_io_rob_commit_0_valid; // @[Core.scala 39:16]
  assign io_rob_commit_0_bits_des_rob = exu_io_rob_commit_0_bits_des_rob; // @[Core.scala 39:16]
  assign io_rob_commit_1_valid = exu_io_rob_commit_1_valid; // @[Core.scala 39:16]
  assign io_rob_commit_1_bits_des_rob = exu_io_rob_commit_1_bits_des_rob; // @[Core.scala 39:16]
  assign io_icache_debug_state = ifu_io_icache_debug_state; // @[Core.scala 42:18]
  assign io_icache_debug_hit_cache = ifu_io_icache_debug_hit_cache; // @[Core.scala 42:18]
  assign io_icache_debug_cache_we = ifu_io_icache_debug_cache_we; // @[Core.scala 42:18]
  assign io_icache_debug_cache_read_tag = ifu_io_icache_debug_cache_read_tag; // @[Core.scala 42:18]
  assign io_icache_debug_icache_req_valid = ifu_io_icache_debug_icache_req_valid; // @[Core.scala 42:18]
  assign io_icache_debug_icache_req_bits_addr = ifu_io_icache_debug_icache_req_bits_addr; // @[Core.scala 42:18]
  assign io_bpu_debug_branch_mask = ifu_io_bpu_debug_branch_mask; // @[Core.scala 43:15]
  assign io_bpu_debug_fetched_mask = ifu_io_bpu_debug_fetched_mask; // @[Core.scala 43:15]
  assign io_bpu_debug_predict_branch = ifu_io_bpu_debug_predict_branch; // @[Core.scala 43:15]
  assign io_bpu_debug_predict_addr = ifu_io_bpu_debug_predict_addr; // @[Core.scala 43:15]
  assign io_bpu_debug_is_taken = ifu_io_bpu_debug_is_taken; // @[Core.scala 43:15]
  assign io_bpu_debug_take_delay = ifu_io_bpu_debug_take_delay; // @[Core.scala 43:15]
  assign io_bpu_debug_inst_packet_0 = ifu_io_bpu_debug_inst_packet_0; // @[Core.scala 43:15]
  assign io_bpu_debug_inst_packet_1 = ifu_io_bpu_debug_inst_packet_1; // @[Core.scala 43:15]
  assign io_bpu_debug_inst_packet_2 = ifu_io_bpu_debug_inst_packet_2; // @[Core.scala 43:15]
  assign io_bpu_debug_inst_packet_3 = ifu_io_bpu_debug_inst_packet_3; // @[Core.scala 43:15]
  assign io_bpu_debug_inst_packet_4 = ifu_io_bpu_debug_inst_packet_4; // @[Core.scala 43:15]
  assign io_bpu_debug_inst_packet_5 = ifu_io_bpu_debug_inst_packet_5; // @[Core.scala 43:15]
  assign io_bpu_debug_inst_packet_6 = ifu_io_bpu_debug_inst_packet_6; // @[Core.scala 43:15]
  assign io_bpu_debug_inst_packet_7 = ifu_io_bpu_debug_inst_packet_7; // @[Core.scala 43:15]
  assign ifu_clock = clock;
  assign ifu_reset = reset;
  assign ifu_io_ex_branch_info_i_valid = exu_io_ex_branch_info_o_valid; // @[Core.scala 29:26]
  assign ifu_io_ex_branch_info_i_bits_target_addr = exu_io_ex_branch_info_o_bits_target_addr; // @[Core.scala 29:26]
  assign ifu_io_ex_branch_info_i_bits_inst_addr = exu_io_ex_branch_info_o_bits_inst_addr; // @[Core.scala 29:26]
  assign ifu_io_ex_branch_info_i_bits_gh_update = exu_io_ex_branch_info_o_bits_gh_update; // @[Core.scala 29:26]
  assign ifu_io_ex_branch_info_i_bits_is_branch = exu_io_ex_branch_info_o_bits_is_branch; // @[Core.scala 29:26]
  assign ifu_io_ex_branch_info_i_bits_is_taken = exu_io_ex_branch_info_o_bits_is_taken; // @[Core.scala 29:26]
  assign ifu_io_ex_branch_info_i_bits_predict_miss = exu_io_ex_branch_info_o_bits_predict_miss; // @[Core.scala 29:26]
  assign ifu_io_fb_resp_deq_valid_0 = exu_io_fb_resp_deq_valid_0; // @[Core.scala 28:17]
  assign ifu_io_fb_resp_deq_valid_1 = exu_io_fb_resp_deq_valid_1; // @[Core.scala 28:17]
  assign ifu_io_icache_io_read_req_ready = io_icache_io_read_req_ready; // @[Core.scala 31:24]
  assign ifu_io_icache_io_read_resp_bits_data = io_icache_io_read_resp_bits_data; // @[Core.scala 32:25]
  assign exu_clock = clock;
  assign exu_reset = reset;
  assign exu_io_fb_inst_bank_i_valid = ifu_io_fb_inst_bank_o_valid; // @[Core.scala 27:24]
  assign exu_io_fb_inst_bank_i_bits_data_0_inst = ifu_io_fb_inst_bank_o_bits_data_0_inst; // @[Core.scala 27:24]
  assign exu_io_fb_inst_bank_i_bits_data_0_inst_addr = ifu_io_fb_inst_bank_o_bits_data_0_inst_addr; // @[Core.scala 27:24]
  assign exu_io_fb_inst_bank_i_bits_data_0_gh_backup = ifu_io_fb_inst_bank_o_bits_data_0_gh_backup; // @[Core.scala 27:24]
  assign exu_io_fb_inst_bank_i_bits_data_0_is_valid = ifu_io_fb_inst_bank_o_bits_data_0_is_valid; // @[Core.scala 27:24]
  assign exu_io_fb_inst_bank_i_bits_data_0_predict_taken = ifu_io_fb_inst_bank_o_bits_data_0_predict_taken; // @[Core.scala 27:24]
  assign exu_io_fb_inst_bank_i_bits_data_1_inst = ifu_io_fb_inst_bank_o_bits_data_1_inst; // @[Core.scala 27:24]
  assign exu_io_fb_inst_bank_i_bits_data_1_inst_addr = ifu_io_fb_inst_bank_o_bits_data_1_inst_addr; // @[Core.scala 27:24]
  assign exu_io_fb_inst_bank_i_bits_data_1_gh_backup = ifu_io_fb_inst_bank_o_bits_data_1_gh_backup; // @[Core.scala 27:24]
  assign exu_io_fb_inst_bank_i_bits_data_1_is_valid = ifu_io_fb_inst_bank_o_bits_data_1_is_valid; // @[Core.scala 27:24]
  assign exu_io_fb_inst_bank_i_bits_data_1_predict_taken = ifu_io_fb_inst_bank_o_bits_data_1_predict_taken; // @[Core.scala 27:24]
  assign exu_io_dcache_io_read_req_ready = io_dcache_io_read_req_ready; // @[Core.scala 34:25]
  assign exu_io_dcache_io_read_resp_bits_data = io_dcache_io_read_resp_bits_data; // @[Core.scala 35:25]
  assign exu_io_dcache_io_write_req_ready = io_dcache_io_write_req_ready; // @[Core.scala 36:25]
endmodule
module IoControl(
  input          clock,
  input          reset,
  output         io_icache_read_req_ready,
  input          io_icache_read_req_valid,
  input  [31:0]  io_icache_read_req_bits_addr,
  output [255:0] io_icache_read_resp_bits_data,
  output         io_dcache_read_req_ready,
  input          io_dcache_read_req_valid,
  input  [31:0]  io_dcache_read_req_bits_addr,
  input  [3:0]   io_dcache_read_req_bits_rob_idx,
  output [31:0]  io_dcache_read_resp_bits_data,
  output         io_dcache_write_req_ready,
  input          io_dcache_write_req_valid,
  input  [31:0]  io_dcache_write_req_bits_addr,
  input  [31:0]  io_dcache_write_req_bits_data,
  input  [3:0]   io_dcache_write_req_bits_byte_mask,
  input  [31:0]  io_base_ram_ctrl_data_in,
  output [31:0]  io_base_ram_ctrl_ctrl_data_out,
  output [19:0]  io_base_ram_ctrl_ctrl_addr,
  output [3:0]   io_base_ram_ctrl_ctrl_be_n,
  output         io_base_ram_ctrl_ctrl_ce_n,
  output         io_base_ram_ctrl_ctrl_oe_n,
  output         io_base_ram_ctrl_ctrl_we_n,
  input  [31:0]  io_ext_ram_ctrl_data_in,
  output [31:0]  io_ext_ram_ctrl_ctrl_data_out,
  output [19:0]  io_ext_ram_ctrl_ctrl_addr,
  output [3:0]   io_ext_ram_ctrl_ctrl_be_n,
  output         io_ext_ram_ctrl_ctrl_ce_n,
  output         io_ext_ram_ctrl_ctrl_oe_n,
  output         io_ext_ram_ctrl_ctrl_we_n,
  input          io_rxd_uart_ready,
  output         io_rxd_uart_clear,
  input  [7:0]   io_rxd_uart_data,
  output         io_txd_uart_start,
  output [7:0]   io_txd_uart_data,
  input          io_txd_uart_busy,
  input          io_rob_commit_0_valid,
  input  [2:0]   io_rob_commit_0_bits_des_rob,
  input          io_rob_commit_1_valid,
  input  [2:0]   io_rob_commit_1_bits_des_rob,
  input          io_need_flush,
  output [2:0]   io_debug_base_state,
  output         io_debug_icache_read_base,
  output         io_debug_icache_read_ext,
  output         io_debug_dcache_read_base,
  output         io_debug_dcache_read_ext,
  output         io_debug_dcache_write_base,
  output         io_debug_dcache_write_ext,
  output [19:0]  io_debug_icache_read_addr,
  output [19:0]  io_debug_dcache_read_addr,
  output [19:0]  io_debug_dcache_write_addr
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [31:0] _RAND_57;
  reg [31:0] _RAND_58;
  reg [31:0] _RAND_59;
  reg [31:0] _RAND_60;
  reg [31:0] _RAND_61;
`endif // RANDOMIZE_REG_INIT
  reg [31:0] base_ram_ctrl_data_out; // @[IoControl.scala 114:26]
  reg [19:0] base_ram_ctrl_addr; // @[IoControl.scala 114:26]
  reg [3:0] base_ram_ctrl_be_n; // @[IoControl.scala 114:26]
  reg  base_ram_ctrl_ce_n; // @[IoControl.scala 114:26]
  reg  base_ram_ctrl_oe_n; // @[IoControl.scala 114:26]
  reg  base_ram_ctrl_we_n; // @[IoControl.scala 114:26]
  reg [31:0] ext_ram_ctrl_data_out; // @[IoControl.scala 115:26]
  reg [19:0] ext_ram_ctrl_addr; // @[IoControl.scala 115:26]
  reg [3:0] ext_ram_ctrl_be_n; // @[IoControl.scala 115:26]
  reg  ext_ram_ctrl_ce_n; // @[IoControl.scala 115:26]
  reg  ext_ram_ctrl_oe_n; // @[IoControl.scala 115:26]
  reg  ext_ram_ctrl_we_n; // @[IoControl.scala 115:26]
  reg [2:0] base_state; // @[IoControl.scala 120:46]
  reg [3:0] base_clock_counter; // @[IoControl.scala 121:46]
  reg [3:0] base_wait_counter; // @[IoControl.scala 122:45]
  reg [2:0] ext_state; // @[IoControl.scala 123:46]
  reg [3:0] ext_clock_counter; // @[IoControl.scala 124:46]
  reg [3:0] ext_wait_counter; // @[IoControl.scala 125:45]
  wire  icache_read_base = io_icache_read_req_bits_addr[31:22] == 10'h200 & io_icache_read_req_valid; // @[IoControl.scala 127:101]
  wire  icache_read_ext = io_icache_read_req_bits_addr[31:22] == 10'h201 & io_icache_read_req_valid; // @[IoControl.scala 128:101]
  wire  dcache_read_base = io_dcache_read_req_bits_addr[31:22] == 10'h200 & io_dcache_read_req_valid; // @[IoControl.scala 129:101]
  wire  dcache_read_ext = io_dcache_read_req_bits_addr[31:22] == 10'h201 & io_dcache_read_req_valid; // @[IoControl.scala 130:101]
  wire  dcache_write_base = io_dcache_write_req_bits_addr[31:22] == 10'h200 & io_dcache_write_req_valid; // @[IoControl.scala 131:102]
  wire  dcache_write_ext = io_dcache_write_req_bits_addr[31:22] == 10'h201 & io_dcache_write_req_valid; // @[IoControl.scala 132:102]
  wire  dcache_read_uart = io_dcache_read_req_bits_addr == 32'hbfd003f8 & io_dcache_read_req_valid; // @[IoControl.scala 133:92]
  wire  dcache_write_uart = io_dcache_write_req_bits_addr == 32'hbfd003f8 & io_dcache_write_req_valid; // @[IoControl.scala 134:94]
  wire  dcache_read_uart_state = io_dcache_read_req_bits_addr == 32'hbfd003fc & io_dcache_read_req_valid; // @[IoControl.scala 135:91]
  wire [19:0] icache_read_addr = io_icache_read_req_bits_addr[21:2]; // @[IoControl.scala 136:67]
  wire [19:0] dcache_read_addr = io_dcache_read_req_bits_addr[21:2]; // @[IoControl.scala 137:67]
  wire [19:0] dcache_write_addr = io_dcache_write_req_bits_addr[21:2]; // @[IoControl.scala 138:68]
  wire  _icache_read_other_T = ~icache_read_base; // @[IoControl.scala 139:27]
  wire  _icache_read_other_T_1 = ~icache_read_ext; // @[IoControl.scala 139:47]
  wire  icache_read_other = ~icache_read_base & ~icache_read_ext & io_icache_read_req_valid; // @[IoControl.scala 139:64]
  wire  _dcache_read_other_T = ~dcache_read_base; // @[IoControl.scala 140:27]
  wire  _dcache_read_other_T_1 = ~dcache_read_ext; // @[IoControl.scala 140:47]
  wire  dcache_read_other = ~dcache_read_base & ~dcache_read_ext & ~dcache_read_uart & io_dcache_read_req_valid; // @[IoControl.scala 140:85]
  wire  _dcache_write_other_T = ~dcache_write_base; // @[IoControl.scala 141:28]
  wire  _dcache_write_other_T_1 = ~dcache_write_ext; // @[IoControl.scala 141:49]
  wire  dcache_write_other = ~dcache_write_base & ~dcache_write_ext & ~dcache_write_uart & io_dcache_write_req_valid; // @[IoControl.scala 141:89]
  reg [31:0] icache_buffer_0; // @[IoControl.scala 155:34]
  reg [31:0] icache_buffer_1; // @[IoControl.scala 155:34]
  reg [31:0] icache_buffer_2; // @[IoControl.scala 155:34]
  reg [31:0] icache_buffer_3; // @[IoControl.scala 155:34]
  reg [31:0] icache_buffer_4; // @[IoControl.scala 155:34]
  reg [31:0] icache_buffer_5; // @[IoControl.scala 155:34]
  reg [31:0] icache_buffer_6; // @[IoControl.scala 155:34]
  reg [31:0] icache_buffer_7; // @[IoControl.scala 155:34]
  reg  icache_data_valid; // @[IoControl.scala 156:34]
  wire [127:0] io_icache_read_resp_bits_data_lo = {icache_buffer_3,icache_buffer_2,icache_buffer_1,icache_buffer_0}; // @[IoControl.scala 159:56]
  wire [127:0] io_icache_read_resp_bits_data_hi = {icache_buffer_7,icache_buffer_6,icache_buffer_5,icache_buffer_4}; // @[IoControl.scala 159:56]
  reg [31:0] dcache_buffer; // @[IoControl.scala 160:34]
  reg  dcache_data_valid; // @[IoControl.scala 161:34]
  reg [1:0] other_state; // @[IoControl.scala 169:28]
  wire  _T = 2'h0 == other_state; // @[Conditional.scala 37:30]
  wire [31:0] _GEN_0 = icache_read_other ? 32'h0 : icache_buffer_0; // @[IoControl.scala 173:30 IoControl.scala 174:22 IoControl.scala 155:34]
  wire [31:0] _GEN_1 = icache_read_other ? 32'h0 : icache_buffer_1; // @[IoControl.scala 173:30 IoControl.scala 174:22 IoControl.scala 155:34]
  wire [31:0] _GEN_2 = icache_read_other ? 32'h0 : icache_buffer_2; // @[IoControl.scala 173:30 IoControl.scala 174:22 IoControl.scala 155:34]
  wire [31:0] _GEN_3 = icache_read_other ? 32'h0 : icache_buffer_3; // @[IoControl.scala 173:30 IoControl.scala 174:22 IoControl.scala 155:34]
  wire [31:0] _GEN_4 = icache_read_other ? 32'h0 : icache_buffer_4; // @[IoControl.scala 173:30 IoControl.scala 174:22 IoControl.scala 155:34]
  wire [31:0] _GEN_5 = icache_read_other ? 32'h0 : icache_buffer_5; // @[IoControl.scala 173:30 IoControl.scala 174:22 IoControl.scala 155:34]
  wire [31:0] _GEN_6 = icache_read_other ? 32'h0 : icache_buffer_6; // @[IoControl.scala 173:30 IoControl.scala 174:22 IoControl.scala 155:34]
  wire [31:0] _GEN_7 = icache_read_other ? 32'h0 : icache_buffer_7; // @[IoControl.scala 173:30 IoControl.scala 174:22 IoControl.scala 155:34]
  wire  _GEN_8 = icache_read_other | icache_data_valid; // @[IoControl.scala 173:30 IoControl.scala 175:26 IoControl.scala 156:34]
  wire [1:0] _GEN_9 = icache_read_other ? 2'h1 : other_state; // @[IoControl.scala 173:30 IoControl.scala 176:20 IoControl.scala 169:28]
  wire [31:0] _GEN_10 = dcache_read_other ? 32'h0 : dcache_buffer; // @[IoControl.scala 178:30 IoControl.scala 179:22 IoControl.scala 160:34]
  wire  _GEN_11 = dcache_read_other | dcache_data_valid; // @[IoControl.scala 178:30 IoControl.scala 180:26 IoControl.scala 161:34]
  wire  _T_1 = 2'h1 == other_state; // @[Conditional.scala 37:30]
  wire  _T_2 = 2'h2 == other_state; // @[Conditional.scala 37:30]
  wire  _T_3 = 2'h3 == other_state; // @[Conditional.scala 37:30]
  wire [1:0] _GEN_15 = _T_3 ? 2'h0 : other_state; // @[Conditional.scala 39:67 IoControl.scala 197:18 IoControl.scala 169:28]
  wire  _GEN_16 = _T_2 ? 1'h0 : dcache_data_valid; // @[Conditional.scala 39:67 IoControl.scala 193:24 IoControl.scala 161:34]
  wire  _GEN_18 = _T_1 ? 1'h0 : icache_data_valid; // @[Conditional.scala 39:67 IoControl.scala 189:24 IoControl.scala 156:34]
  wire  _GEN_20 = _T_1 ? dcache_data_valid : _GEN_16; // @[Conditional.scala 39:67 IoControl.scala 161:34]
  wire [31:0] _GEN_21 = _T ? _GEN_0 : icache_buffer_0; // @[Conditional.scala 40:58 IoControl.scala 155:34]
  wire [31:0] _GEN_22 = _T ? _GEN_1 : icache_buffer_1; // @[Conditional.scala 40:58 IoControl.scala 155:34]
  wire [31:0] _GEN_23 = _T ? _GEN_2 : icache_buffer_2; // @[Conditional.scala 40:58 IoControl.scala 155:34]
  wire [31:0] _GEN_24 = _T ? _GEN_3 : icache_buffer_3; // @[Conditional.scala 40:58 IoControl.scala 155:34]
  wire [31:0] _GEN_25 = _T ? _GEN_4 : icache_buffer_4; // @[Conditional.scala 40:58 IoControl.scala 155:34]
  wire [31:0] _GEN_26 = _T ? _GEN_5 : icache_buffer_5; // @[Conditional.scala 40:58 IoControl.scala 155:34]
  wire [31:0] _GEN_27 = _T ? _GEN_6 : icache_buffer_6; // @[Conditional.scala 40:58 IoControl.scala 155:34]
  wire [31:0] _GEN_28 = _T ? _GEN_7 : icache_buffer_7; // @[Conditional.scala 40:58 IoControl.scala 155:34]
  wire  _GEN_29 = _T ? _GEN_8 : _GEN_18; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_31 = _T ? _GEN_10 : dcache_buffer; // @[Conditional.scala 40:58 IoControl.scala 160:34]
  wire  _GEN_32 = _T ? _GEN_11 : _GEN_20; // @[Conditional.scala 40:58]
  wire  _GEN_33 = _T & dcache_write_other; // @[Conditional.scala 40:58]
  wire  _T_4 = 3'h0 == base_state; // @[Conditional.scala 37:30]
  wire [3:0] _T_5 = ~io_dcache_write_req_bits_byte_mask; // @[IoControl.scala 209:129]
  wire [2:0] _GEN_34 = icache_read_base ? 3'h1 : base_state; // @[IoControl.scala 217:36 IoControl.scala 218:20 IoControl.scala 120:46]
  wire [31:0] _GEN_35 = icache_read_base ? 32'h0 : base_ram_ctrl_data_out; // @[IoControl.scala 217:36 IoControl.scala 21:14 IoControl.scala 114:26]
  wire [19:0] _GEN_36 = icache_read_base ? icache_read_addr : base_ram_ctrl_addr; // @[IoControl.scala 217:36 IoControl.scala 22:10 IoControl.scala 114:26]
  wire [3:0] _GEN_37 = icache_read_base ? 4'h0 : base_ram_ctrl_be_n; // @[IoControl.scala 217:36 IoControl.scala 23:10 IoControl.scala 114:26]
  wire  _GEN_38 = icache_read_base ? 1'h0 : base_ram_ctrl_ce_n; // @[IoControl.scala 217:36 IoControl.scala 24:10 IoControl.scala 114:26]
  wire  _GEN_39 = icache_read_base ? 1'h0 : base_ram_ctrl_oe_n; // @[IoControl.scala 217:36 IoControl.scala 25:10 IoControl.scala 114:26]
  wire  _GEN_40 = icache_read_base | base_ram_ctrl_we_n; // @[IoControl.scala 217:36 IoControl.scala 26:10 IoControl.scala 114:26]
  wire [3:0] _GEN_41 = icache_read_base ? 4'h0 : base_clock_counter; // @[IoControl.scala 217:36 IoControl.scala 220:28 IoControl.scala 121:46]
  wire [3:0] _GEN_42 = icache_read_base ? 4'h0 : base_wait_counter; // @[IoControl.scala 217:36 IoControl.scala 221:27 IoControl.scala 122:45]
  wire  _GEN_47 = dcache_read_base ? 1'h0 : _GEN_38; // @[IoControl.scala 212:36 IoControl.scala 24:10]
  wire  _GEN_48 = dcache_read_base ? 1'h0 : _GEN_39; // @[IoControl.scala 212:36 IoControl.scala 25:10]
  wire  _GEN_49 = dcache_read_base | _GEN_40; // @[IoControl.scala 212:36 IoControl.scala 26:10]
  wire  _GEN_56 = dcache_write_base ? 1'h0 : _GEN_47; // @[IoControl.scala 206:31 IoControl.scala 33:10]
  wire  _GEN_57 = dcache_write_base | _GEN_48; // @[IoControl.scala 206:31 IoControl.scala 34:10]
  wire  _GEN_58 = dcache_write_base ? 1'h0 : _GEN_49; // @[IoControl.scala 206:31 IoControl.scala 35:10]
  wire  _T_6 = 3'h1 == base_state; // @[Conditional.scala 37:30]
  wire  _T_9 = base_wait_counter == 4'h1; // @[IoControl.scala 231:32]
  wire [31:0] _GEN_61 = 3'h0 == base_clock_counter[2:0] ? io_base_ram_ctrl_data_in : _GEN_21; // @[IoControl.scala 232:45 IoControl.scala 232:45]
  wire [31:0] _GEN_62 = 3'h1 == base_clock_counter[2:0] ? io_base_ram_ctrl_data_in : _GEN_22; // @[IoControl.scala 232:45 IoControl.scala 232:45]
  wire [31:0] _GEN_63 = 3'h2 == base_clock_counter[2:0] ? io_base_ram_ctrl_data_in : _GEN_23; // @[IoControl.scala 232:45 IoControl.scala 232:45]
  wire [31:0] _GEN_64 = 3'h3 == base_clock_counter[2:0] ? io_base_ram_ctrl_data_in : _GEN_24; // @[IoControl.scala 232:45 IoControl.scala 232:45]
  wire [31:0] _GEN_65 = 3'h4 == base_clock_counter[2:0] ? io_base_ram_ctrl_data_in : _GEN_25; // @[IoControl.scala 232:45 IoControl.scala 232:45]
  wire [31:0] _GEN_66 = 3'h5 == base_clock_counter[2:0] ? io_base_ram_ctrl_data_in : _GEN_26; // @[IoControl.scala 232:45 IoControl.scala 232:45]
  wire [31:0] _GEN_67 = 3'h6 == base_clock_counter[2:0] ? io_base_ram_ctrl_data_in : _GEN_27; // @[IoControl.scala 232:45 IoControl.scala 232:45]
  wire [31:0] _GEN_68 = 3'h7 == base_clock_counter[2:0] ? io_base_ram_ctrl_data_in : _GEN_28; // @[IoControl.scala 232:45 IoControl.scala 232:45]
  wire [3:0] _base_wait_counter_T_1 = base_wait_counter + 4'h1; // @[IoControl.scala 238:47]
  wire [31:0] _GEN_69 = base_wait_counter == 4'h1 ? _GEN_61 : _GEN_21; // @[IoControl.scala 231:49]
  wire [31:0] _GEN_70 = base_wait_counter == 4'h1 ? _GEN_62 : _GEN_22; // @[IoControl.scala 231:49]
  wire [31:0] _GEN_71 = base_wait_counter == 4'h1 ? _GEN_63 : _GEN_23; // @[IoControl.scala 231:49]
  wire [31:0] _GEN_72 = base_wait_counter == 4'h1 ? _GEN_64 : _GEN_24; // @[IoControl.scala 231:49]
  wire [31:0] _GEN_73 = base_wait_counter == 4'h1 ? _GEN_65 : _GEN_25; // @[IoControl.scala 231:49]
  wire [31:0] _GEN_74 = base_wait_counter == 4'h1 ? _GEN_66 : _GEN_26; // @[IoControl.scala 231:49]
  wire [31:0] _GEN_75 = base_wait_counter == 4'h1 ? _GEN_67 : _GEN_27; // @[IoControl.scala 231:49]
  wire [31:0] _GEN_76 = base_wait_counter == 4'h1 ? _GEN_68 : _GEN_28; // @[IoControl.scala 231:49]
  wire [31:0] _GEN_77 = base_wait_counter == 4'h1 ? 32'h0 : base_ram_ctrl_data_out; // @[IoControl.scala 231:49 IoControl.scala 12:14 IoControl.scala 114:26]
  wire [19:0] _GEN_78 = base_wait_counter == 4'h1 ? 20'h0 : base_ram_ctrl_addr; // @[IoControl.scala 231:49 IoControl.scala 13:10 IoControl.scala 114:26]
  wire [3:0] _GEN_79 = base_wait_counter == 4'h1 ? 4'hf : base_ram_ctrl_be_n; // @[IoControl.scala 231:49 IoControl.scala 14:10 IoControl.scala 114:26]
  wire  _GEN_80 = base_wait_counter == 4'h1 | base_ram_ctrl_ce_n; // @[IoControl.scala 231:49 IoControl.scala 15:10 IoControl.scala 114:26]
  wire  _GEN_81 = base_wait_counter == 4'h1 | base_ram_ctrl_oe_n; // @[IoControl.scala 231:49 IoControl.scala 16:10 IoControl.scala 114:26]
  wire  _GEN_82 = base_wait_counter == 4'h1 | base_ram_ctrl_we_n; // @[IoControl.scala 231:49 IoControl.scala 17:10 IoControl.scala 114:26]
  wire  _GEN_83 = base_wait_counter == 4'h1 | _GEN_29; // @[IoControl.scala 231:49 IoControl.scala 234:29]
  wire [2:0] _GEN_84 = base_wait_counter == 4'h1 ? 3'h4 : base_state; // @[IoControl.scala 231:49 IoControl.scala 235:22 IoControl.scala 120:46]
  wire [3:0] _GEN_85 = base_wait_counter == 4'h1 ? 4'h0 : _base_wait_counter_T_1; // @[IoControl.scala 231:49 IoControl.scala 236:28 IoControl.scala 238:28]
  wire [19:0] _T_13 = base_ram_ctrl_addr + 20'h1; // @[IoControl.scala 242:49]
  wire [3:0] _base_clock_counter_T_1 = base_clock_counter + 4'h1; // @[IoControl.scala 244:52]
  wire [19:0] _GEN_95 = _T_9 ? _T_13 : base_ram_ctrl_addr; // @[IoControl.scala 241:48 IoControl.scala 22:10 IoControl.scala 114:26]
  wire [3:0] _GEN_96 = _T_9 ? 4'h0 : base_ram_ctrl_be_n; // @[IoControl.scala 241:48 IoControl.scala 23:10 IoControl.scala 114:26]
  wire  _GEN_97 = _T_9 ? 1'h0 : base_ram_ctrl_ce_n; // @[IoControl.scala 241:48 IoControl.scala 24:10 IoControl.scala 114:26]
  wire  _GEN_98 = _T_9 ? 1'h0 : base_ram_ctrl_oe_n; // @[IoControl.scala 241:48 IoControl.scala 25:10 IoControl.scala 114:26]
  wire [3:0] _GEN_108 = _T_9 ? _base_clock_counter_T_1 : base_clock_counter; // @[IoControl.scala 241:48 IoControl.scala 244:30 IoControl.scala 121:46]
  wire [31:0] _GEN_110 = base_clock_counter == 4'h7 ? _GEN_69 : _GEN_69; // @[IoControl.scala 230:60]
  wire [31:0] _GEN_111 = base_clock_counter == 4'h7 ? _GEN_70 : _GEN_70; // @[IoControl.scala 230:60]
  wire [31:0] _GEN_112 = base_clock_counter == 4'h7 ? _GEN_71 : _GEN_71; // @[IoControl.scala 230:60]
  wire [31:0] _GEN_113 = base_clock_counter == 4'h7 ? _GEN_72 : _GEN_72; // @[IoControl.scala 230:60]
  wire [31:0] _GEN_114 = base_clock_counter == 4'h7 ? _GEN_73 : _GEN_73; // @[IoControl.scala 230:60]
  wire [31:0] _GEN_115 = base_clock_counter == 4'h7 ? _GEN_74 : _GEN_74; // @[IoControl.scala 230:60]
  wire [31:0] _GEN_116 = base_clock_counter == 4'h7 ? _GEN_75 : _GEN_75; // @[IoControl.scala 230:60]
  wire [31:0] _GEN_117 = base_clock_counter == 4'h7 ? _GEN_76 : _GEN_76; // @[IoControl.scala 230:60]
  wire [31:0] _GEN_118 = base_clock_counter == 4'h7 ? _GEN_77 : _GEN_77; // @[IoControl.scala 230:60]
  wire [19:0] _GEN_119 = base_clock_counter == 4'h7 ? _GEN_78 : _GEN_95; // @[IoControl.scala 230:60]
  wire [3:0] _GEN_120 = base_clock_counter == 4'h7 ? _GEN_79 : _GEN_96; // @[IoControl.scala 230:60]
  wire  _GEN_121 = base_clock_counter == 4'h7 ? _GEN_80 : _GEN_97; // @[IoControl.scala 230:60]
  wire  _GEN_122 = base_clock_counter == 4'h7 ? _GEN_81 : _GEN_98; // @[IoControl.scala 230:60]
  wire  _GEN_123 = base_clock_counter == 4'h7 ? _GEN_82 : _GEN_82; // @[IoControl.scala 230:60]
  wire  _GEN_124 = base_clock_counter == 4'h7 ? _GEN_83 : _GEN_29; // @[IoControl.scala 230:60]
  wire [2:0] _GEN_125 = base_clock_counter == 4'h7 ? _GEN_84 : base_state; // @[IoControl.scala 230:60 IoControl.scala 120:46]
  wire [3:0] _GEN_126 = base_clock_counter == 4'h7 ? _GEN_85 : _GEN_85; // @[IoControl.scala 230:60]
  wire [3:0] _GEN_127 = base_clock_counter == 4'h7 ? base_clock_counter : _GEN_108; // @[IoControl.scala 230:60 IoControl.scala 121:46]
  wire  _GEN_131 = _icache_read_other_T | _GEN_121; // @[IoControl.scala 225:31 IoControl.scala 15:10]
  wire  _GEN_132 = _icache_read_other_T | _GEN_122; // @[IoControl.scala 225:31 IoControl.scala 16:10]
  wire  _GEN_133 = _icache_read_other_T | _GEN_123; // @[IoControl.scala 225:31 IoControl.scala 17:10]
  wire [31:0] _GEN_137 = _icache_read_other_T ? _GEN_21 : _GEN_110; // @[IoControl.scala 225:31]
  wire [31:0] _GEN_138 = _icache_read_other_T ? _GEN_22 : _GEN_111; // @[IoControl.scala 225:31]
  wire [31:0] _GEN_139 = _icache_read_other_T ? _GEN_23 : _GEN_112; // @[IoControl.scala 225:31]
  wire [31:0] _GEN_140 = _icache_read_other_T ? _GEN_24 : _GEN_113; // @[IoControl.scala 225:31]
  wire [31:0] _GEN_141 = _icache_read_other_T ? _GEN_25 : _GEN_114; // @[IoControl.scala 225:31]
  wire [31:0] _GEN_142 = _icache_read_other_T ? _GEN_26 : _GEN_115; // @[IoControl.scala 225:31]
  wire [31:0] _GEN_143 = _icache_read_other_T ? _GEN_27 : _GEN_116; // @[IoControl.scala 225:31]
  wire [31:0] _GEN_144 = _icache_read_other_T ? _GEN_28 : _GEN_117; // @[IoControl.scala 225:31]
  wire  _GEN_145 = _icache_read_other_T ? _GEN_29 : _GEN_124; // @[IoControl.scala 225:31]
  wire  _T_15 = 3'h4 == base_state; // @[Conditional.scala 37:30]
  wire  _T_16 = 3'h2 == base_state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_146 = _T_9 ? 3'h5 : base_state; // @[IoControl.scala 261:52 IoControl.scala 262:20 IoControl.scala 120:46]
  wire [31:0] _GEN_153 = _T_9 ? io_base_ram_ctrl_data_in : _GEN_31; // @[IoControl.scala 261:52 IoControl.scala 264:23]
  wire  _GEN_154 = _T_9 | _GEN_32; // @[IoControl.scala 261:52 IoControl.scala 265:27]
  wire [3:0] _GEN_155 = _T_9 ? base_wait_counter : _base_wait_counter_T_1; // @[IoControl.scala 261:52 IoControl.scala 122:45 IoControl.scala 267:26]
  wire [31:0] _GEN_156 = _dcache_read_other_T ? 32'h0 : _GEN_77; // @[IoControl.scala 256:31 IoControl.scala 12:14]
  wire [19:0] _GEN_157 = _dcache_read_other_T ? 20'h0 : _GEN_78; // @[IoControl.scala 256:31 IoControl.scala 13:10]
  wire [3:0] _GEN_158 = _dcache_read_other_T ? 4'hf : _GEN_79; // @[IoControl.scala 256:31 IoControl.scala 14:10]
  wire  _GEN_159 = _dcache_read_other_T | _GEN_80; // @[IoControl.scala 256:31 IoControl.scala 15:10]
  wire  _GEN_160 = _dcache_read_other_T | _GEN_81; // @[IoControl.scala 256:31 IoControl.scala 16:10]
  wire  _GEN_161 = _dcache_read_other_T | _GEN_82; // @[IoControl.scala 256:31 IoControl.scala 17:10]
  wire [2:0] _GEN_162 = _dcache_read_other_T ? 3'h0 : _GEN_146; // @[IoControl.scala 256:31 IoControl.scala 258:20]
  wire [3:0] _GEN_163 = _dcache_read_other_T ? 4'h0 : base_clock_counter; // @[IoControl.scala 256:31 IoControl.scala 259:28 IoControl.scala 121:46]
  wire [3:0] _GEN_164 = _dcache_read_other_T ? 4'h0 : _GEN_155; // @[IoControl.scala 256:31 IoControl.scala 260:27]
  wire [31:0] _GEN_165 = _dcache_read_other_T ? _GEN_31 : _GEN_153; // @[IoControl.scala 256:31]
  wire  _GEN_166 = _dcache_read_other_T ? _GEN_32 : _GEN_154; // @[IoControl.scala 256:31]
  wire  _T_19 = 3'h5 == base_state; // @[Conditional.scala 37:30]
  wire  _T_20 = 3'h3 == base_state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_167 = _T_9 ? 3'h0 : base_state; // @[IoControl.scala 280:52 IoControl.scala 281:20 IoControl.scala 120:46]
  wire  _GEN_174 = _T_9 | _GEN_33; // @[IoControl.scala 280:52 IoControl.scala 283:31]
  wire [31:0] _GEN_176 = _dcache_write_other_T ? 32'h0 : _GEN_77; // @[IoControl.scala 275:32 IoControl.scala 12:14]
  wire [19:0] _GEN_177 = _dcache_write_other_T ? 20'h0 : _GEN_78; // @[IoControl.scala 275:32 IoControl.scala 13:10]
  wire [3:0] _GEN_178 = _dcache_write_other_T ? 4'hf : _GEN_79; // @[IoControl.scala 275:32 IoControl.scala 14:10]
  wire  _GEN_179 = _dcache_write_other_T | _GEN_80; // @[IoControl.scala 275:32 IoControl.scala 15:10]
  wire  _GEN_180 = _dcache_write_other_T | _GEN_81; // @[IoControl.scala 275:32 IoControl.scala 16:10]
  wire  _GEN_181 = _dcache_write_other_T | _GEN_82; // @[IoControl.scala 275:32 IoControl.scala 17:10]
  wire [2:0] _GEN_182 = _dcache_write_other_T ? 3'h0 : _GEN_167; // @[IoControl.scala 275:32 IoControl.scala 277:20]
  wire [3:0] _GEN_183 = _dcache_write_other_T ? 4'h0 : base_clock_counter; // @[IoControl.scala 275:32 IoControl.scala 278:28 IoControl.scala 121:46]
  wire [3:0] _GEN_184 = _dcache_write_other_T ? 4'h0 : _GEN_155; // @[IoControl.scala 275:32 IoControl.scala 279:27]
  wire  _GEN_185 = _dcache_write_other_T ? _GEN_33 : _GEN_174; // @[IoControl.scala 275:32]
  wire [31:0] _GEN_186 = _T_20 ? _GEN_176 : base_ram_ctrl_data_out; // @[Conditional.scala 39:67 IoControl.scala 114:26]
  wire [19:0] _GEN_187 = _T_20 ? _GEN_177 : base_ram_ctrl_addr; // @[Conditional.scala 39:67 IoControl.scala 114:26]
  wire [3:0] _GEN_188 = _T_20 ? _GEN_178 : base_ram_ctrl_be_n; // @[Conditional.scala 39:67 IoControl.scala 114:26]
  wire  _GEN_189 = _T_20 ? _GEN_179 : base_ram_ctrl_ce_n; // @[Conditional.scala 39:67 IoControl.scala 114:26]
  wire  _GEN_190 = _T_20 ? _GEN_180 : base_ram_ctrl_oe_n; // @[Conditional.scala 39:67 IoControl.scala 114:26]
  wire  _GEN_191 = _T_20 ? _GEN_181 : base_ram_ctrl_we_n; // @[Conditional.scala 39:67 IoControl.scala 114:26]
  wire [2:0] _GEN_192 = _T_20 ? _GEN_182 : base_state; // @[Conditional.scala 39:67 IoControl.scala 120:46]
  wire [3:0] _GEN_193 = _T_20 ? _GEN_183 : base_clock_counter; // @[Conditional.scala 39:67 IoControl.scala 121:46]
  wire [3:0] _GEN_194 = _T_20 ? _GEN_184 : base_wait_counter; // @[Conditional.scala 39:67 IoControl.scala 122:45]
  wire  _GEN_195 = _T_20 ? _GEN_185 : _GEN_33; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_196 = _T_19 ? 3'h0 : _GEN_192; // @[Conditional.scala 39:67 IoControl.scala 271:20]
  wire  _GEN_197 = _T_19 ? 1'h0 : _GEN_32; // @[Conditional.scala 39:67 IoControl.scala 272:27]
  wire [31:0] _GEN_198 = _T_19 ? base_ram_ctrl_data_out : _GEN_186; // @[Conditional.scala 39:67 IoControl.scala 114:26]
  wire [19:0] _GEN_199 = _T_19 ? base_ram_ctrl_addr : _GEN_187; // @[Conditional.scala 39:67 IoControl.scala 114:26]
  wire [3:0] _GEN_200 = _T_19 ? base_ram_ctrl_be_n : _GEN_188; // @[Conditional.scala 39:67 IoControl.scala 114:26]
  wire  _GEN_201 = _T_19 ? base_ram_ctrl_ce_n : _GEN_189; // @[Conditional.scala 39:67 IoControl.scala 114:26]
  wire  _GEN_202 = _T_19 ? base_ram_ctrl_oe_n : _GEN_190; // @[Conditional.scala 39:67 IoControl.scala 114:26]
  wire  _GEN_203 = _T_19 ? base_ram_ctrl_we_n : _GEN_191; // @[Conditional.scala 39:67 IoControl.scala 114:26]
  wire [3:0] _GEN_204 = _T_19 ? base_clock_counter : _GEN_193; // @[Conditional.scala 39:67 IoControl.scala 121:46]
  wire [3:0] _GEN_205 = _T_19 ? base_wait_counter : _GEN_194; // @[Conditional.scala 39:67 IoControl.scala 122:45]
  wire  _GEN_206 = _T_19 ? _GEN_33 : _GEN_195; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_207 = _T_16 ? _GEN_156 : _GEN_198; // @[Conditional.scala 39:67]
  wire [19:0] _GEN_208 = _T_16 ? _GEN_157 : _GEN_199; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_209 = _T_16 ? _GEN_158 : _GEN_200; // @[Conditional.scala 39:67]
  wire  _GEN_210 = _T_16 ? _GEN_159 : _GEN_201; // @[Conditional.scala 39:67]
  wire  _GEN_211 = _T_16 ? _GEN_160 : _GEN_202; // @[Conditional.scala 39:67]
  wire  _GEN_212 = _T_16 ? _GEN_161 : _GEN_203; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_213 = _T_16 ? _GEN_162 : _GEN_196; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_214 = _T_16 ? _GEN_163 : _GEN_204; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_215 = _T_16 ? _GEN_164 : _GEN_205; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_216 = _T_16 ? _GEN_165 : _GEN_31; // @[Conditional.scala 39:67]
  wire  _GEN_217 = _T_16 ? _GEN_166 : _GEN_197; // @[Conditional.scala 39:67]
  wire  _GEN_218 = _T_16 ? _GEN_33 : _GEN_206; // @[Conditional.scala 39:67]
  wire  _GEN_220 = _T_15 ? 1'h0 : _GEN_29; // @[Conditional.scala 39:67 IoControl.scala 253:27]
  wire  _GEN_224 = _T_15 ? base_ram_ctrl_ce_n : _GEN_210; // @[Conditional.scala 39:67 IoControl.scala 114:26]
  wire  _GEN_225 = _T_15 ? base_ram_ctrl_oe_n : _GEN_211; // @[Conditional.scala 39:67 IoControl.scala 114:26]
  wire  _GEN_226 = _T_15 ? base_ram_ctrl_we_n : _GEN_212; // @[Conditional.scala 39:67 IoControl.scala 114:26]
  wire [31:0] _GEN_229 = _T_15 ? _GEN_31 : _GEN_216; // @[Conditional.scala 39:67]
  wire  _GEN_230 = _T_15 ? _GEN_32 : _GEN_217; // @[Conditional.scala 39:67]
  wire  _GEN_231 = _T_15 ? _GEN_33 : _GEN_218; // @[Conditional.scala 39:67]
  wire  _GEN_235 = _T_6 ? _GEN_131 : _GEN_224; // @[Conditional.scala 39:67]
  wire  _GEN_236 = _T_6 ? _GEN_132 : _GEN_225; // @[Conditional.scala 39:67]
  wire  _GEN_237 = _T_6 ? _GEN_133 : _GEN_226; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_241 = _T_6 ? _GEN_137 : _GEN_21; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_242 = _T_6 ? _GEN_138 : _GEN_22; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_243 = _T_6 ? _GEN_139 : _GEN_23; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_244 = _T_6 ? _GEN_140 : _GEN_24; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_245 = _T_6 ? _GEN_141 : _GEN_25; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_246 = _T_6 ? _GEN_142 : _GEN_26; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_247 = _T_6 ? _GEN_143 : _GEN_27; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_248 = _T_6 ? _GEN_144 : _GEN_28; // @[Conditional.scala 39:67]
  wire  _GEN_249 = _T_6 ? _GEN_145 : _GEN_220; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_250 = _T_6 ? _GEN_31 : _GEN_229; // @[Conditional.scala 39:67]
  wire  _GEN_251 = _T_6 ? _GEN_32 : _GEN_230; // @[Conditional.scala 39:67]
  wire  _GEN_252 = _T_6 ? _GEN_33 : _GEN_231; // @[Conditional.scala 39:67]
  wire  _GEN_257 = _T_4 ? _GEN_56 : _GEN_235; // @[Conditional.scala 40:58]
  wire  _GEN_258 = _T_4 ? _GEN_57 : _GEN_236; // @[Conditional.scala 40:58]
  wire  _GEN_259 = _T_4 ? _GEN_58 : _GEN_237; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_262 = _T_4 ? _GEN_21 : _GEN_241; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_263 = _T_4 ? _GEN_22 : _GEN_242; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_264 = _T_4 ? _GEN_23 : _GEN_243; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_265 = _T_4 ? _GEN_24 : _GEN_244; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_266 = _T_4 ? _GEN_25 : _GEN_245; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_267 = _T_4 ? _GEN_26 : _GEN_246; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_268 = _T_4 ? _GEN_27 : _GEN_247; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_269 = _T_4 ? _GEN_28 : _GEN_248; // @[Conditional.scala 40:58]
  wire  _GEN_270 = _T_4 ? _GEN_29 : _GEN_249; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_271 = _T_4 ? _GEN_31 : _GEN_250; // @[Conditional.scala 40:58]
  wire  _GEN_272 = _T_4 ? _GEN_32 : _GEN_251; // @[Conditional.scala 40:58]
  wire  _GEN_273 = _T_4 ? _T & dcache_write_other : _GEN_252; // @[Conditional.scala 40:58]
  wire  _T_23 = 3'h0 == ext_state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_274 = icache_read_ext ? 3'h1 : ext_state; // @[IoControl.scala 303:35 IoControl.scala 304:19 IoControl.scala 123:46]
  wire [31:0] _GEN_275 = icache_read_ext ? 32'h0 : ext_ram_ctrl_data_out; // @[IoControl.scala 303:35 IoControl.scala 21:14 IoControl.scala 115:26]
  wire [19:0] _GEN_276 = icache_read_ext ? icache_read_addr : ext_ram_ctrl_addr; // @[IoControl.scala 303:35 IoControl.scala 22:10 IoControl.scala 115:26]
  wire [3:0] _GEN_277 = icache_read_ext ? 4'h0 : ext_ram_ctrl_be_n; // @[IoControl.scala 303:35 IoControl.scala 23:10 IoControl.scala 115:26]
  wire  _GEN_278 = icache_read_ext ? 1'h0 : ext_ram_ctrl_ce_n; // @[IoControl.scala 303:35 IoControl.scala 24:10 IoControl.scala 115:26]
  wire  _GEN_279 = icache_read_ext ? 1'h0 : ext_ram_ctrl_oe_n; // @[IoControl.scala 303:35 IoControl.scala 25:10 IoControl.scala 115:26]
  wire  _GEN_280 = icache_read_ext | ext_ram_ctrl_we_n; // @[IoControl.scala 303:35 IoControl.scala 26:10 IoControl.scala 115:26]
  wire [3:0] _GEN_281 = icache_read_ext ? 4'h0 : ext_clock_counter; // @[IoControl.scala 303:35 IoControl.scala 306:27 IoControl.scala 124:46]
  wire [3:0] _GEN_282 = icache_read_ext ? 4'h0 : ext_wait_counter; // @[IoControl.scala 303:35 IoControl.scala 307:26 IoControl.scala 125:45]
  wire  _GEN_287 = dcache_write_ext ? 1'h0 : _GEN_278; // @[IoControl.scala 297:36 IoControl.scala 33:10]
  wire  _GEN_288 = dcache_write_ext | _GEN_279; // @[IoControl.scala 297:36 IoControl.scala 34:10]
  wire  _GEN_289 = dcache_write_ext ? 1'h0 : _GEN_280; // @[IoControl.scala 297:36 IoControl.scala 35:10]
  wire  _GEN_296 = dcache_read_ext ? 1'h0 : _GEN_287; // @[IoControl.scala 292:29 IoControl.scala 24:10]
  wire  _GEN_297 = dcache_read_ext ? 1'h0 : _GEN_288; // @[IoControl.scala 292:29 IoControl.scala 25:10]
  wire  _GEN_298 = dcache_read_ext | _GEN_289; // @[IoControl.scala 292:29 IoControl.scala 26:10]
  wire  _T_25 = 3'h1 == ext_state; // @[Conditional.scala 37:30]
  wire  _T_28 = ext_wait_counter == 4'h1; // @[IoControl.scala 317:31]
  wire [31:0] _GEN_301 = 3'h0 == ext_clock_counter[2:0] ? io_ext_ram_ctrl_data_in : _GEN_262; // @[IoControl.scala 318:44 IoControl.scala 318:44]
  wire [31:0] _GEN_302 = 3'h1 == ext_clock_counter[2:0] ? io_ext_ram_ctrl_data_in : _GEN_263; // @[IoControl.scala 318:44 IoControl.scala 318:44]
  wire [31:0] _GEN_303 = 3'h2 == ext_clock_counter[2:0] ? io_ext_ram_ctrl_data_in : _GEN_264; // @[IoControl.scala 318:44 IoControl.scala 318:44]
  wire [31:0] _GEN_304 = 3'h3 == ext_clock_counter[2:0] ? io_ext_ram_ctrl_data_in : _GEN_265; // @[IoControl.scala 318:44 IoControl.scala 318:44]
  wire [31:0] _GEN_305 = 3'h4 == ext_clock_counter[2:0] ? io_ext_ram_ctrl_data_in : _GEN_266; // @[IoControl.scala 318:44 IoControl.scala 318:44]
  wire [31:0] _GEN_306 = 3'h5 == ext_clock_counter[2:0] ? io_ext_ram_ctrl_data_in : _GEN_267; // @[IoControl.scala 318:44 IoControl.scala 318:44]
  wire [31:0] _GEN_307 = 3'h6 == ext_clock_counter[2:0] ? io_ext_ram_ctrl_data_in : _GEN_268; // @[IoControl.scala 318:44 IoControl.scala 318:44]
  wire [31:0] _GEN_308 = 3'h7 == ext_clock_counter[2:0] ? io_ext_ram_ctrl_data_in : _GEN_269; // @[IoControl.scala 318:44 IoControl.scala 318:44]
  wire [3:0] _ext_wait_counter_T_1 = ext_wait_counter + 4'h1; // @[IoControl.scala 324:45]
  wire [31:0] _GEN_309 = ext_wait_counter == 4'h1 ? _GEN_301 : _GEN_262; // @[IoControl.scala 317:47]
  wire [31:0] _GEN_310 = ext_wait_counter == 4'h1 ? _GEN_302 : _GEN_263; // @[IoControl.scala 317:47]
  wire [31:0] _GEN_311 = ext_wait_counter == 4'h1 ? _GEN_303 : _GEN_264; // @[IoControl.scala 317:47]
  wire [31:0] _GEN_312 = ext_wait_counter == 4'h1 ? _GEN_304 : _GEN_265; // @[IoControl.scala 317:47]
  wire [31:0] _GEN_313 = ext_wait_counter == 4'h1 ? _GEN_305 : _GEN_266; // @[IoControl.scala 317:47]
  wire [31:0] _GEN_314 = ext_wait_counter == 4'h1 ? _GEN_306 : _GEN_267; // @[IoControl.scala 317:47]
  wire [31:0] _GEN_315 = ext_wait_counter == 4'h1 ? _GEN_307 : _GEN_268; // @[IoControl.scala 317:47]
  wire [31:0] _GEN_316 = ext_wait_counter == 4'h1 ? _GEN_308 : _GEN_269; // @[IoControl.scala 317:47]
  wire [31:0] _GEN_317 = ext_wait_counter == 4'h1 ? 32'h0 : ext_ram_ctrl_data_out; // @[IoControl.scala 317:47 IoControl.scala 12:14 IoControl.scala 115:26]
  wire [19:0] _GEN_318 = ext_wait_counter == 4'h1 ? 20'h0 : ext_ram_ctrl_addr; // @[IoControl.scala 317:47 IoControl.scala 13:10 IoControl.scala 115:26]
  wire [3:0] _GEN_319 = ext_wait_counter == 4'h1 ? 4'hf : ext_ram_ctrl_be_n; // @[IoControl.scala 317:47 IoControl.scala 14:10 IoControl.scala 115:26]
  wire  _GEN_320 = ext_wait_counter == 4'h1 | ext_ram_ctrl_ce_n; // @[IoControl.scala 317:47 IoControl.scala 15:10 IoControl.scala 115:26]
  wire  _GEN_321 = ext_wait_counter == 4'h1 | ext_ram_ctrl_oe_n; // @[IoControl.scala 317:47 IoControl.scala 16:10 IoControl.scala 115:26]
  wire  _GEN_322 = ext_wait_counter == 4'h1 | ext_ram_ctrl_we_n; // @[IoControl.scala 317:47 IoControl.scala 17:10 IoControl.scala 115:26]
  wire  _GEN_323 = ext_wait_counter == 4'h1 | _GEN_270; // @[IoControl.scala 317:47 IoControl.scala 320:29]
  wire [2:0] _GEN_324 = ext_wait_counter == 4'h1 ? 3'h4 : ext_state; // @[IoControl.scala 317:47 IoControl.scala 321:21 IoControl.scala 123:46]
  wire [3:0] _GEN_325 = ext_wait_counter == 4'h1 ? 4'h0 : _ext_wait_counter_T_1; // @[IoControl.scala 317:47 IoControl.scala 322:27 IoControl.scala 324:27]
  wire [19:0] _T_32 = ext_ram_ctrl_addr + 20'h1; // @[IoControl.scala 328:47]
  wire [3:0] _ext_clock_counter_T_1 = ext_clock_counter + 4'h1; // @[IoControl.scala 330:50]
  wire [19:0] _GEN_335 = _T_28 ? _T_32 : ext_ram_ctrl_addr; // @[IoControl.scala 327:47 IoControl.scala 22:10 IoControl.scala 115:26]
  wire [3:0] _GEN_336 = _T_28 ? 4'h0 : ext_ram_ctrl_be_n; // @[IoControl.scala 327:47 IoControl.scala 23:10 IoControl.scala 115:26]
  wire  _GEN_337 = _T_28 ? 1'h0 : ext_ram_ctrl_ce_n; // @[IoControl.scala 327:47 IoControl.scala 24:10 IoControl.scala 115:26]
  wire  _GEN_338 = _T_28 ? 1'h0 : ext_ram_ctrl_oe_n; // @[IoControl.scala 327:47 IoControl.scala 25:10 IoControl.scala 115:26]
  wire [3:0] _GEN_348 = _T_28 ? _ext_clock_counter_T_1 : ext_clock_counter; // @[IoControl.scala 327:47 IoControl.scala 330:29 IoControl.scala 124:46]
  wire [31:0] _GEN_350 = ext_clock_counter == 4'h7 ? _GEN_309 : _GEN_309; // @[IoControl.scala 316:59]
  wire [31:0] _GEN_351 = ext_clock_counter == 4'h7 ? _GEN_310 : _GEN_310; // @[IoControl.scala 316:59]
  wire [31:0] _GEN_352 = ext_clock_counter == 4'h7 ? _GEN_311 : _GEN_311; // @[IoControl.scala 316:59]
  wire [31:0] _GEN_353 = ext_clock_counter == 4'h7 ? _GEN_312 : _GEN_312; // @[IoControl.scala 316:59]
  wire [31:0] _GEN_354 = ext_clock_counter == 4'h7 ? _GEN_313 : _GEN_313; // @[IoControl.scala 316:59]
  wire [31:0] _GEN_355 = ext_clock_counter == 4'h7 ? _GEN_314 : _GEN_314; // @[IoControl.scala 316:59]
  wire [31:0] _GEN_356 = ext_clock_counter == 4'h7 ? _GEN_315 : _GEN_315; // @[IoControl.scala 316:59]
  wire [31:0] _GEN_357 = ext_clock_counter == 4'h7 ? _GEN_316 : _GEN_316; // @[IoControl.scala 316:59]
  wire [31:0] _GEN_358 = ext_clock_counter == 4'h7 ? _GEN_317 : _GEN_317; // @[IoControl.scala 316:59]
  wire [19:0] _GEN_359 = ext_clock_counter == 4'h7 ? _GEN_318 : _GEN_335; // @[IoControl.scala 316:59]
  wire [3:0] _GEN_360 = ext_clock_counter == 4'h7 ? _GEN_319 : _GEN_336; // @[IoControl.scala 316:59]
  wire  _GEN_361 = ext_clock_counter == 4'h7 ? _GEN_320 : _GEN_337; // @[IoControl.scala 316:59]
  wire  _GEN_362 = ext_clock_counter == 4'h7 ? _GEN_321 : _GEN_338; // @[IoControl.scala 316:59]
  wire  _GEN_363 = ext_clock_counter == 4'h7 ? _GEN_322 : _GEN_322; // @[IoControl.scala 316:59]
  wire  _GEN_364 = ext_clock_counter == 4'h7 ? _GEN_323 : _GEN_270; // @[IoControl.scala 316:59]
  wire [2:0] _GEN_365 = ext_clock_counter == 4'h7 ? _GEN_324 : ext_state; // @[IoControl.scala 316:59 IoControl.scala 123:46]
  wire [3:0] _GEN_366 = ext_clock_counter == 4'h7 ? _GEN_325 : _GEN_325; // @[IoControl.scala 316:59]
  wire [3:0] _GEN_367 = ext_clock_counter == 4'h7 ? ext_clock_counter : _GEN_348; // @[IoControl.scala 316:59 IoControl.scala 124:46]
  wire  _GEN_371 = _icache_read_other_T_1 | _GEN_361; // @[IoControl.scala 311:30 IoControl.scala 15:10]
  wire  _GEN_372 = _icache_read_other_T_1 | _GEN_362; // @[IoControl.scala 311:30 IoControl.scala 16:10]
  wire  _GEN_373 = _icache_read_other_T_1 | _GEN_363; // @[IoControl.scala 311:30 IoControl.scala 17:10]
  wire  _T_34 = 3'h4 == ext_state; // @[Conditional.scala 37:30]
  wire  _T_35 = 3'h2 == ext_state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_386 = _T_28 ? 3'h5 : ext_state; // @[IoControl.scala 347:51 IoControl.scala 348:19 IoControl.scala 123:46]
  wire [31:0] _GEN_393 = _T_28 ? io_ext_ram_ctrl_data_in : _GEN_271; // @[IoControl.scala 347:51 IoControl.scala 350:23]
  wire  _GEN_394 = _T_28 | _GEN_272; // @[IoControl.scala 347:51 IoControl.scala 351:27]
  wire [3:0] _GEN_395 = _T_28 ? ext_wait_counter : _ext_wait_counter_T_1; // @[IoControl.scala 347:51 IoControl.scala 125:45 IoControl.scala 353:25]
  wire [31:0] _GEN_396 = _dcache_read_other_T_1 ? 32'h0 : _GEN_317; // @[IoControl.scala 342:30 IoControl.scala 12:14]
  wire [19:0] _GEN_397 = _dcache_read_other_T_1 ? 20'h0 : _GEN_318; // @[IoControl.scala 342:30 IoControl.scala 13:10]
  wire [3:0] _GEN_398 = _dcache_read_other_T_1 ? 4'hf : _GEN_319; // @[IoControl.scala 342:30 IoControl.scala 14:10]
  wire  _GEN_399 = _dcache_read_other_T_1 | _GEN_320; // @[IoControl.scala 342:30 IoControl.scala 15:10]
  wire  _GEN_400 = _dcache_read_other_T_1 | _GEN_321; // @[IoControl.scala 342:30 IoControl.scala 16:10]
  wire  _GEN_401 = _dcache_read_other_T_1 | _GEN_322; // @[IoControl.scala 342:30 IoControl.scala 17:10]
  wire [2:0] _GEN_402 = _dcache_read_other_T_1 ? 3'h0 : _GEN_386; // @[IoControl.scala 342:30 IoControl.scala 344:19]
  wire [3:0] _GEN_403 = _dcache_read_other_T_1 ? 4'h0 : ext_clock_counter; // @[IoControl.scala 342:30 IoControl.scala 345:27 IoControl.scala 124:46]
  wire [3:0] _GEN_404 = _dcache_read_other_T_1 ? 4'h0 : _GEN_395; // @[IoControl.scala 342:30 IoControl.scala 346:26]
  wire [31:0] _GEN_405 = _dcache_read_other_T_1 ? _GEN_271 : _GEN_393; // @[IoControl.scala 342:30]
  wire  _GEN_406 = _dcache_read_other_T_1 ? _GEN_272 : _GEN_394; // @[IoControl.scala 342:30]
  wire  _T_38 = 3'h5 == ext_state; // @[Conditional.scala 37:30]
  wire  _T_39 = 3'h3 == ext_state; // @[Conditional.scala 37:30]
  wire [2:0] _GEN_407 = _T_28 ? 3'h0 : ext_state; // @[IoControl.scala 366:51 IoControl.scala 367:19 IoControl.scala 123:46]
  wire  _GEN_414 = _T_28 | _GEN_273; // @[IoControl.scala 366:51 IoControl.scala 369:31]
  wire [31:0] _GEN_416 = _dcache_write_other_T_1 ? 32'h0 : _GEN_317; // @[IoControl.scala 361:31 IoControl.scala 12:14]
  wire [19:0] _GEN_417 = _dcache_write_other_T_1 ? 20'h0 : _GEN_318; // @[IoControl.scala 361:31 IoControl.scala 13:10]
  wire [3:0] _GEN_418 = _dcache_write_other_T_1 ? 4'hf : _GEN_319; // @[IoControl.scala 361:31 IoControl.scala 14:10]
  wire  _GEN_419 = _dcache_write_other_T_1 | _GEN_320; // @[IoControl.scala 361:31 IoControl.scala 15:10]
  wire  _GEN_420 = _dcache_write_other_T_1 | _GEN_321; // @[IoControl.scala 361:31 IoControl.scala 16:10]
  wire  _GEN_421 = _dcache_write_other_T_1 | _GEN_322; // @[IoControl.scala 361:31 IoControl.scala 17:10]
  wire [2:0] _GEN_422 = _dcache_write_other_T_1 ? 3'h0 : _GEN_407; // @[IoControl.scala 361:31 IoControl.scala 363:19]
  wire [3:0] _GEN_423 = _dcache_write_other_T_1 ? 4'h0 : ext_clock_counter; // @[IoControl.scala 361:31 IoControl.scala 364:27 IoControl.scala 124:46]
  wire [3:0] _GEN_424 = _dcache_write_other_T_1 ? 4'h0 : _GEN_395; // @[IoControl.scala 361:31 IoControl.scala 365:26]
  wire  _GEN_425 = _dcache_write_other_T_1 ? _GEN_273 : _GEN_414; // @[IoControl.scala 361:31]
  wire [31:0] _GEN_426 = _T_39 ? _GEN_416 : ext_ram_ctrl_data_out; // @[Conditional.scala 39:67 IoControl.scala 115:26]
  wire [19:0] _GEN_427 = _T_39 ? _GEN_417 : ext_ram_ctrl_addr; // @[Conditional.scala 39:67 IoControl.scala 115:26]
  wire [3:0] _GEN_428 = _T_39 ? _GEN_418 : ext_ram_ctrl_be_n; // @[Conditional.scala 39:67 IoControl.scala 115:26]
  wire  _GEN_429 = _T_39 ? _GEN_419 : ext_ram_ctrl_ce_n; // @[Conditional.scala 39:67 IoControl.scala 115:26]
  wire  _GEN_430 = _T_39 ? _GEN_420 : ext_ram_ctrl_oe_n; // @[Conditional.scala 39:67 IoControl.scala 115:26]
  wire  _GEN_431 = _T_39 ? _GEN_421 : ext_ram_ctrl_we_n; // @[Conditional.scala 39:67 IoControl.scala 115:26]
  wire [2:0] _GEN_432 = _T_39 ? _GEN_422 : ext_state; // @[Conditional.scala 39:67 IoControl.scala 123:46]
  wire [3:0] _GEN_433 = _T_39 ? _GEN_423 : ext_clock_counter; // @[Conditional.scala 39:67 IoControl.scala 124:46]
  wire [3:0] _GEN_434 = _T_39 ? _GEN_424 : ext_wait_counter; // @[Conditional.scala 39:67 IoControl.scala 125:45]
  wire  _GEN_435 = _T_39 ? _GEN_425 : _GEN_273; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_436 = _T_38 ? 3'h0 : _GEN_432; // @[Conditional.scala 39:67 IoControl.scala 357:17]
  wire  _GEN_437 = _T_38 ? 1'h0 : _GEN_272; // @[Conditional.scala 39:67 IoControl.scala 358:25]
  wire [31:0] _GEN_438 = _T_38 ? ext_ram_ctrl_data_out : _GEN_426; // @[Conditional.scala 39:67 IoControl.scala 115:26]
  wire [19:0] _GEN_439 = _T_38 ? ext_ram_ctrl_addr : _GEN_427; // @[Conditional.scala 39:67 IoControl.scala 115:26]
  wire [3:0] _GEN_440 = _T_38 ? ext_ram_ctrl_be_n : _GEN_428; // @[Conditional.scala 39:67 IoControl.scala 115:26]
  wire  _GEN_441 = _T_38 ? ext_ram_ctrl_ce_n : _GEN_429; // @[Conditional.scala 39:67 IoControl.scala 115:26]
  wire  _GEN_442 = _T_38 ? ext_ram_ctrl_oe_n : _GEN_430; // @[Conditional.scala 39:67 IoControl.scala 115:26]
  wire  _GEN_443 = _T_38 ? ext_ram_ctrl_we_n : _GEN_431; // @[Conditional.scala 39:67 IoControl.scala 115:26]
  wire [3:0] _GEN_444 = _T_38 ? ext_clock_counter : _GEN_433; // @[Conditional.scala 39:67 IoControl.scala 124:46]
  wire [3:0] _GEN_445 = _T_38 ? ext_wait_counter : _GEN_434; // @[Conditional.scala 39:67 IoControl.scala 125:45]
  wire  _GEN_446 = _T_38 ? _GEN_273 : _GEN_435; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_447 = _T_35 ? _GEN_396 : _GEN_438; // @[Conditional.scala 39:67]
  wire [19:0] _GEN_448 = _T_35 ? _GEN_397 : _GEN_439; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_449 = _T_35 ? _GEN_398 : _GEN_440; // @[Conditional.scala 39:67]
  wire  _GEN_450 = _T_35 ? _GEN_399 : _GEN_441; // @[Conditional.scala 39:67]
  wire  _GEN_451 = _T_35 ? _GEN_400 : _GEN_442; // @[Conditional.scala 39:67]
  wire  _GEN_452 = _T_35 ? _GEN_401 : _GEN_443; // @[Conditional.scala 39:67]
  wire [2:0] _GEN_453 = _T_35 ? _GEN_402 : _GEN_436; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_454 = _T_35 ? _GEN_403 : _GEN_444; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_455 = _T_35 ? _GEN_404 : _GEN_445; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_456 = _T_35 ? _GEN_405 : _GEN_271; // @[Conditional.scala 39:67]
  wire  _GEN_457 = _T_35 ? _GEN_406 : _GEN_437; // @[Conditional.scala 39:67]
  wire  _GEN_458 = _T_35 ? _GEN_273 : _GEN_446; // @[Conditional.scala 39:67]
  wire  _GEN_464 = _T_34 ? ext_ram_ctrl_ce_n : _GEN_450; // @[Conditional.scala 39:67 IoControl.scala 115:26]
  wire  _GEN_465 = _T_34 ? ext_ram_ctrl_oe_n : _GEN_451; // @[Conditional.scala 39:67 IoControl.scala 115:26]
  wire  _GEN_466 = _T_34 ? ext_ram_ctrl_we_n : _GEN_452; // @[Conditional.scala 39:67 IoControl.scala 115:26]
  wire [31:0] _GEN_469 = _T_34 ? _GEN_271 : _GEN_456; // @[Conditional.scala 39:67]
  wire  _GEN_470 = _T_34 ? _GEN_272 : _GEN_457; // @[Conditional.scala 39:67]
  wire  _GEN_471 = _T_34 ? _GEN_273 : _GEN_458; // @[Conditional.scala 39:67]
  wire  _GEN_475 = _T_25 ? _GEN_371 : _GEN_464; // @[Conditional.scala 39:67]
  wire  _GEN_476 = _T_25 ? _GEN_372 : _GEN_465; // @[Conditional.scala 39:67]
  wire  _GEN_477 = _T_25 ? _GEN_373 : _GEN_466; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_490 = _T_25 ? _GEN_271 : _GEN_469; // @[Conditional.scala 39:67]
  wire  _GEN_491 = _T_25 ? _GEN_272 : _GEN_470; // @[Conditional.scala 39:67]
  wire  _GEN_492 = _T_25 ? _GEN_273 : _GEN_471; // @[Conditional.scala 39:67]
  wire  _GEN_497 = _T_23 ? _GEN_296 : _GEN_475; // @[Conditional.scala 40:58]
  wire  _GEN_498 = _T_23 ? _GEN_297 : _GEN_476; // @[Conditional.scala 40:58]
  wire  _GEN_499 = _T_23 ? _GEN_298 : _GEN_477; // @[Conditional.scala 40:58]
  wire [31:0] _GEN_511 = _T_23 ? _GEN_271 : _GEN_490; // @[Conditional.scala 40:58]
  wire  _GEN_512 = _T_23 ? _GEN_272 : _GEN_491; // @[Conditional.scala 40:58]
  wire  _GEN_513 = _T_23 ? _GEN_273 : _GEN_492; // @[Conditional.scala 40:58]
  reg [7:0] uart_buffer_0_data; // @[IoControl.scala 378:24]
  reg [2:0] uart_buffer_0_rob_idx; // @[IoControl.scala 378:24]
  reg [7:0] uart_buffer_1_data; // @[IoControl.scala 378:24]
  reg [2:0] uart_buffer_1_rob_idx; // @[IoControl.scala 378:24]
  reg [7:0] uart_buffer_2_data; // @[IoControl.scala 378:24]
  reg [2:0] uart_buffer_2_rob_idx; // @[IoControl.scala 378:24]
  reg [7:0] uart_buffer_3_data; // @[IoControl.scala 378:24]
  reg [2:0] uart_buffer_3_rob_idx; // @[IoControl.scala 378:24]
  reg [7:0] uart_buffer_4_data; // @[IoControl.scala 378:24]
  reg [2:0] uart_buffer_4_rob_idx; // @[IoControl.scala 378:24]
  reg [7:0] uart_buffer_5_data; // @[IoControl.scala 378:24]
  reg [2:0] uart_buffer_5_rob_idx; // @[IoControl.scala 378:24]
  reg [7:0] uart_buffer_6_data; // @[IoControl.scala 378:24]
  reg [2:0] uart_buffer_6_rob_idx; // @[IoControl.scala 378:24]
  reg [7:0] uart_buffer_7_data; // @[IoControl.scala 378:24]
  reg [2:0] uart_buffer_7_rob_idx; // @[IoControl.scala 378:24]
  reg  uart_buffer_wait_0; // @[IoControl.scala 379:33]
  reg  uart_buffer_wait_1; // @[IoControl.scala 379:33]
  reg  uart_buffer_wait_2; // @[IoControl.scala 379:33]
  reg  uart_buffer_wait_3; // @[IoControl.scala 379:33]
  reg  uart_buffer_wait_4; // @[IoControl.scala 379:33]
  reg  uart_buffer_wait_5; // @[IoControl.scala 379:33]
  reg  uart_buffer_wait_6; // @[IoControl.scala 379:33]
  reg  uart_buffer_wait_7; // @[IoControl.scala 379:33]
  reg [7:0] uart_head; // @[IoControl.scala 380:26]
  wire [3:0] head_idx_hi = uart_head[7:4]; // @[OneHot.scala 30:18]
  wire [3:0] head_idx_lo = uart_head[3:0]; // @[OneHot.scala 31:18]
  wire  head_idx_hi_1 = |head_idx_hi; // @[OneHot.scala 32:14]
  wire [3:0] _head_idx_T = head_idx_hi | head_idx_lo; // @[OneHot.scala 32:28]
  wire [1:0] head_idx_hi_2 = _head_idx_T[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] head_idx_lo_1 = _head_idx_T[1:0]; // @[OneHot.scala 31:18]
  wire  head_idx_hi_3 = |head_idx_hi_2; // @[OneHot.scala 32:14]
  wire [1:0] _head_idx_T_1 = head_idx_hi_2 | head_idx_lo_1; // @[OneHot.scala 32:28]
  wire  head_idx_lo_2 = _head_idx_T_1[1]; // @[CircuitMath.scala 30:8]
  wire [2:0] head_idx = {head_idx_hi_1,head_idx_hi_3,head_idx_lo_2}; // @[Cat.scala 30:58]
  reg [7:0] uart_flush_head; // @[IoControl.scala 382:32]
  reg [7:0] uart_tail; // @[IoControl.scala 383:26]
  wire [3:0] tail_idx_hi = uart_tail[7:4]; // @[OneHot.scala 30:18]
  wire [3:0] tail_idx_lo = uart_tail[3:0]; // @[OneHot.scala 31:18]
  wire  tail_idx_hi_1 = |tail_idx_hi; // @[OneHot.scala 32:14]
  wire [3:0] _tail_idx_T = tail_idx_hi | tail_idx_lo; // @[OneHot.scala 32:28]
  wire [1:0] tail_idx_hi_2 = _tail_idx_T[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] tail_idx_lo_1 = _tail_idx_T[1:0]; // @[OneHot.scala 31:18]
  wire  tail_idx_hi_3 = |tail_idx_hi_2; // @[OneHot.scala 32:14]
  wire [1:0] _tail_idx_T_1 = tail_idx_hi_2 | tail_idx_lo_1; // @[OneHot.scala 32:28]
  wire  tail_idx_lo_2 = _tail_idx_T_1[1]; // @[CircuitMath.scala 30:8]
  wire [2:0] tail_idx = {tail_idx_hi_1,tail_idx_hi_3,tail_idx_lo_2}; // @[Cat.scala 30:58]
  reg  maybe_full; // @[IoControl.scala 385:27]
  reg  maybe_true_full; // @[IoControl.scala 386:32]
  wire  uart_full = uart_flush_head == uart_tail & maybe_true_full; // @[IoControl.scala 387:46]
  wire  uart_empty = uart_head == uart_tail & ~maybe_full; // @[IoControl.scala 388:41]
  wire  _uart_enq_T = ~uart_full; // @[IoControl.scala 396:18]
  wire  write_req = io_rxd_uart_ready & _uart_enq_T; // @[IoControl.scala 458:25]
  wire  uart_enq = ~uart_full & write_req; // @[IoControl.scala 396:28]
  wire  _uart_deq_T = ~uart_empty; // @[IoControl.scala 397:18]
  reg [1:0] uart_state; // @[IoControl.scala 452:27]
  wire  _T_56 = 2'h0 == uart_state; // @[Conditional.scala 37:30]
  wire  _T_57 = ~io_txd_uart_busy; // @[IoControl.scala 470:32]
  wire  _T_59 = dcache_read_uart & _uart_deq_T; // @[IoControl.scala 475:34]
  wire  _GEN_782 = dcache_write_uart & ~io_txd_uart_busy ? 1'h0 : _T_59; // @[IoControl.scala 470:50]
  wire  read_req = _T_56 & _GEN_782; // @[Conditional.scala 40:58]
  wire  uart_deq = ~uart_empty & read_req; // @[IoControl.scala 397:29]
  wire [7:0] _GEN_515 = 3'h1 == head_idx ? uart_buffer_1_data : uart_buffer_0_data; // @[IoControl.scala 399:12 IoControl.scala 399:12]
  wire [7:0] _GEN_516 = 3'h2 == head_idx ? uart_buffer_2_data : _GEN_515; // @[IoControl.scala 399:12 IoControl.scala 399:12]
  wire [7:0] _GEN_517 = 3'h3 == head_idx ? uart_buffer_3_data : _GEN_516; // @[IoControl.scala 399:12 IoControl.scala 399:12]
  wire [7:0] _GEN_518 = 3'h4 == head_idx ? uart_buffer_4_data : _GEN_517; // @[IoControl.scala 399:12 IoControl.scala 399:12]
  wire [7:0] _GEN_519 = 3'h5 == head_idx ? uart_buffer_5_data : _GEN_518; // @[IoControl.scala 399:12 IoControl.scala 399:12]
  wire [7:0] _GEN_520 = 3'h6 == head_idx ? uart_buffer_6_data : _GEN_519; // @[IoControl.scala 399:12 IoControl.scala 399:12]
  wire [7:0] read_data = 3'h7 == head_idx ? uart_buffer_7_data : _GEN_520; // @[IoControl.scala 399:12 IoControl.scala 399:12]
  wire [2:0] _GEN_530 = 3'h0 == tail_idx ? 3'h0 : uart_buffer_0_rob_idx; // @[IoControl.scala 405:34 IoControl.scala 405:34 IoControl.scala 378:24]
  wire [2:0] _GEN_531 = 3'h1 == tail_idx ? 3'h0 : uart_buffer_1_rob_idx; // @[IoControl.scala 405:34 IoControl.scala 405:34 IoControl.scala 378:24]
  wire [2:0] _GEN_532 = 3'h2 == tail_idx ? 3'h0 : uart_buffer_2_rob_idx; // @[IoControl.scala 405:34 IoControl.scala 405:34 IoControl.scala 378:24]
  wire [2:0] _GEN_533 = 3'h3 == tail_idx ? 3'h0 : uart_buffer_3_rob_idx; // @[IoControl.scala 405:34 IoControl.scala 405:34 IoControl.scala 378:24]
  wire [2:0] _GEN_534 = 3'h4 == tail_idx ? 3'h0 : uart_buffer_4_rob_idx; // @[IoControl.scala 405:34 IoControl.scala 405:34 IoControl.scala 378:24]
  wire [2:0] _GEN_535 = 3'h5 == tail_idx ? 3'h0 : uart_buffer_5_rob_idx; // @[IoControl.scala 405:34 IoControl.scala 405:34 IoControl.scala 378:24]
  wire [2:0] _GEN_536 = 3'h6 == tail_idx ? 3'h0 : uart_buffer_6_rob_idx; // @[IoControl.scala 405:34 IoControl.scala 405:34 IoControl.scala 378:24]
  wire [2:0] _GEN_537 = 3'h7 == tail_idx ? 3'h0 : uart_buffer_7_rob_idx; // @[IoControl.scala 405:34 IoControl.scala 405:34 IoControl.scala 378:24]
  wire [6:0] uart_tail_hi = uart_tail[6:0]; // @[IoControl.scala 106:12]
  wire  uart_tail_lo = uart_tail[7]; // @[IoControl.scala 106:29]
  wire [7:0] _uart_tail_T = {uart_tail_hi,uart_tail_lo}; // @[Cat.scala 30:58]
  wire [2:0] _GEN_546 = uart_enq ? _GEN_530 : uart_buffer_0_rob_idx; // @[IoControl.scala 403:17 IoControl.scala 378:24]
  wire [2:0] _GEN_547 = uart_enq ? _GEN_531 : uart_buffer_1_rob_idx; // @[IoControl.scala 403:17 IoControl.scala 378:24]
  wire [2:0] _GEN_548 = uart_enq ? _GEN_532 : uart_buffer_2_rob_idx; // @[IoControl.scala 403:17 IoControl.scala 378:24]
  wire [2:0] _GEN_549 = uart_enq ? _GEN_533 : uart_buffer_3_rob_idx; // @[IoControl.scala 403:17 IoControl.scala 378:24]
  wire [2:0] _GEN_550 = uart_enq ? _GEN_534 : uart_buffer_4_rob_idx; // @[IoControl.scala 403:17 IoControl.scala 378:24]
  wire [2:0] _GEN_551 = uart_enq ? _GEN_535 : uart_buffer_5_rob_idx; // @[IoControl.scala 403:17 IoControl.scala 378:24]
  wire [2:0] _GEN_552 = uart_enq ? _GEN_536 : uart_buffer_6_rob_idx; // @[IoControl.scala 403:17 IoControl.scala 378:24]
  wire [2:0] _GEN_553 = uart_enq ? _GEN_537 : uart_buffer_7_rob_idx; // @[IoControl.scala 403:17 IoControl.scala 378:24]
  wire [3:0] _GEN_774 = dcache_read_uart & _uart_deq_T ? io_dcache_read_req_bits_rob_idx : 4'h0; // @[IoControl.scala 475:48 IoControl.scala 479:21]
  wire [3:0] _GEN_783 = dcache_write_uart & ~io_txd_uart_busy ? 4'h0 : _GEN_774; // @[IoControl.scala 470:50]
  wire [3:0] _GEN_796 = _T_56 ? _GEN_783 : 4'h0; // @[Conditional.scala 40:58]
  wire [2:0] read_rob_idx = _GEN_796[2:0];
  wire [2:0] _GEN_555 = 3'h0 == head_idx ? read_rob_idx : _GEN_546; // @[IoControl.scala 410:34 IoControl.scala 410:34]
  wire [2:0] _GEN_556 = 3'h1 == head_idx ? read_rob_idx : _GEN_547; // @[IoControl.scala 410:34 IoControl.scala 410:34]
  wire [2:0] _GEN_557 = 3'h2 == head_idx ? read_rob_idx : _GEN_548; // @[IoControl.scala 410:34 IoControl.scala 410:34]
  wire [2:0] _GEN_558 = 3'h3 == head_idx ? read_rob_idx : _GEN_549; // @[IoControl.scala 410:34 IoControl.scala 410:34]
  wire [2:0] _GEN_559 = 3'h4 == head_idx ? read_rob_idx : _GEN_550; // @[IoControl.scala 410:34 IoControl.scala 410:34]
  wire [2:0] _GEN_560 = 3'h5 == head_idx ? read_rob_idx : _GEN_551; // @[IoControl.scala 410:34 IoControl.scala 410:34]
  wire [2:0] _GEN_561 = 3'h6 == head_idx ? read_rob_idx : _GEN_552; // @[IoControl.scala 410:34 IoControl.scala 410:34]
  wire [2:0] _GEN_562 = 3'h7 == head_idx ? read_rob_idx : _GEN_553; // @[IoControl.scala 410:34 IoControl.scala 410:34]
  wire  _GEN_563 = 3'h0 == head_idx | uart_buffer_wait_0; // @[IoControl.scala 411:31 IoControl.scala 411:31 IoControl.scala 379:33]
  wire  _GEN_564 = 3'h1 == head_idx | uart_buffer_wait_1; // @[IoControl.scala 411:31 IoControl.scala 411:31 IoControl.scala 379:33]
  wire  _GEN_565 = 3'h2 == head_idx | uart_buffer_wait_2; // @[IoControl.scala 411:31 IoControl.scala 411:31 IoControl.scala 379:33]
  wire  _GEN_566 = 3'h3 == head_idx | uart_buffer_wait_3; // @[IoControl.scala 411:31 IoControl.scala 411:31 IoControl.scala 379:33]
  wire  _GEN_567 = 3'h4 == head_idx | uart_buffer_wait_4; // @[IoControl.scala 411:31 IoControl.scala 411:31 IoControl.scala 379:33]
  wire  _GEN_568 = 3'h5 == head_idx | uart_buffer_wait_5; // @[IoControl.scala 411:31 IoControl.scala 411:31 IoControl.scala 379:33]
  wire  _GEN_569 = 3'h6 == head_idx | uart_buffer_wait_6; // @[IoControl.scala 411:31 IoControl.scala 411:31 IoControl.scala 379:33]
  wire  _GEN_570 = 3'h7 == head_idx | uart_buffer_wait_7; // @[IoControl.scala 411:31 IoControl.scala 411:31 IoControl.scala 379:33]
  wire [6:0] uart_head_hi = uart_head[6:0]; // @[IoControl.scala 106:12]
  wire  uart_head_lo = uart_head[7]; // @[IoControl.scala 106:29]
  wire [7:0] _uart_head_T = {uart_head_hi,uart_head_lo}; // @[Cat.scala 30:58]
  wire [2:0] _GEN_571 = uart_deq ? _GEN_555 : _GEN_546; // @[IoControl.scala 409:18]
  wire [2:0] _GEN_572 = uart_deq ? _GEN_556 : _GEN_547; // @[IoControl.scala 409:18]
  wire [2:0] _GEN_573 = uart_deq ? _GEN_557 : _GEN_548; // @[IoControl.scala 409:18]
  wire [2:0] _GEN_574 = uart_deq ? _GEN_558 : _GEN_549; // @[IoControl.scala 409:18]
  wire [2:0] _GEN_575 = uart_deq ? _GEN_559 : _GEN_550; // @[IoControl.scala 409:18]
  wire [2:0] _GEN_576 = uart_deq ? _GEN_560 : _GEN_551; // @[IoControl.scala 409:18]
  wire [2:0] _GEN_577 = uart_deq ? _GEN_561 : _GEN_552; // @[IoControl.scala 409:18]
  wire [2:0] _GEN_578 = uart_deq ? _GEN_562 : _GEN_553; // @[IoControl.scala 409:18]
  wire  _GEN_579 = uart_deq ? _GEN_563 : uart_buffer_wait_0; // @[IoControl.scala 409:18 IoControl.scala 379:33]
  wire  _GEN_580 = uart_deq ? _GEN_564 : uart_buffer_wait_1; // @[IoControl.scala 409:18 IoControl.scala 379:33]
  wire  _GEN_581 = uart_deq ? _GEN_565 : uart_buffer_wait_2; // @[IoControl.scala 409:18 IoControl.scala 379:33]
  wire  _GEN_582 = uart_deq ? _GEN_566 : uart_buffer_wait_3; // @[IoControl.scala 409:18 IoControl.scala 379:33]
  wire  _GEN_583 = uart_deq ? _GEN_567 : uart_buffer_wait_4; // @[IoControl.scala 409:18 IoControl.scala 379:33]
  wire  _GEN_584 = uart_deq ? _GEN_568 : uart_buffer_wait_5; // @[IoControl.scala 409:18 IoControl.scala 379:33]
  wire  _GEN_585 = uart_deq ? _GEN_569 : uart_buffer_wait_6; // @[IoControl.scala 409:18 IoControl.scala 379:33]
  wire  _GEN_586 = uart_deq ? _GEN_570 : uart_buffer_wait_7; // @[IoControl.scala 409:18 IoControl.scala 379:33]
  wire [3:0] flush_head_idx_hi = uart_flush_head[7:4]; // @[OneHot.scala 30:18]
  wire [3:0] flush_head_idx_lo = uart_flush_head[3:0]; // @[OneHot.scala 31:18]
  wire  flush_head_idx_hi_1 = |flush_head_idx_hi; // @[OneHot.scala 32:14]
  wire [3:0] _flush_head_idx_T = flush_head_idx_hi | flush_head_idx_lo; // @[OneHot.scala 32:28]
  wire [1:0] flush_head_idx_hi_2 = _flush_head_idx_T[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] flush_head_idx_lo_1 = _flush_head_idx_T[1:0]; // @[OneHot.scala 31:18]
  wire  flush_head_idx_hi_3 = |flush_head_idx_hi_2; // @[OneHot.scala 32:14]
  wire [1:0] _flush_head_idx_T_1 = flush_head_idx_hi_2 | flush_head_idx_lo_1; // @[OneHot.scala 32:28]
  wire  flush_head_idx_lo_2 = _flush_head_idx_T_1[1]; // @[CircuitMath.scala 30:8]
  wire [2:0] flush_head_idx = {flush_head_idx_hi_1,flush_head_idx_hi_3,flush_head_idx_lo_2}; // @[Cat.scala 30:58]
  wire [2:0] _GEN_589 = 3'h1 == flush_head_idx ? uart_buffer_1_rob_idx : uart_buffer_0_rob_idx; // @[IoControl.scala 420:47 IoControl.scala 420:47]
  wire [2:0] _GEN_590 = 3'h2 == flush_head_idx ? uart_buffer_2_rob_idx : _GEN_589; // @[IoControl.scala 420:47 IoControl.scala 420:47]
  wire [2:0] _GEN_591 = 3'h3 == flush_head_idx ? uart_buffer_3_rob_idx : _GEN_590; // @[IoControl.scala 420:47 IoControl.scala 420:47]
  wire [2:0] _GEN_592 = 3'h4 == flush_head_idx ? uart_buffer_4_rob_idx : _GEN_591; // @[IoControl.scala 420:47 IoControl.scala 420:47]
  wire [2:0] _GEN_593 = 3'h5 == flush_head_idx ? uart_buffer_5_rob_idx : _GEN_592; // @[IoControl.scala 420:47 IoControl.scala 420:47]
  wire [2:0] _GEN_594 = 3'h6 == flush_head_idx ? uart_buffer_6_rob_idx : _GEN_593; // @[IoControl.scala 420:47 IoControl.scala 420:47]
  wire [2:0] _GEN_595 = 3'h7 == flush_head_idx ? uart_buffer_7_rob_idx : _GEN_594; // @[IoControl.scala 420:47 IoControl.scala 420:47]
  wire  _GEN_597 = 3'h1 == flush_head_idx ? uart_buffer_wait_1 : uart_buffer_wait_0; // @[IoControl.scala 420:103 IoControl.scala 420:103]
  wire  _GEN_598 = 3'h2 == flush_head_idx ? uart_buffer_wait_2 : _GEN_597; // @[IoControl.scala 420:103 IoControl.scala 420:103]
  wire  _GEN_599 = 3'h3 == flush_head_idx ? uart_buffer_wait_3 : _GEN_598; // @[IoControl.scala 420:103 IoControl.scala 420:103]
  wire  _GEN_600 = 3'h4 == flush_head_idx ? uart_buffer_wait_4 : _GEN_599; // @[IoControl.scala 420:103 IoControl.scala 420:103]
  wire  _GEN_601 = 3'h5 == flush_head_idx ? uart_buffer_wait_5 : _GEN_600; // @[IoControl.scala 420:103 IoControl.scala 420:103]
  wire  _GEN_602 = 3'h6 == flush_head_idx ? uart_buffer_wait_6 : _GEN_601; // @[IoControl.scala 420:103 IoControl.scala 420:103]
  wire  _GEN_603 = 3'h7 == flush_head_idx ? uart_buffer_wait_7 : _GEN_602; // @[IoControl.scala 420:103 IoControl.scala 420:103]
  wire [2:0] _GEN_604 = 3'h0 == flush_head_idx ? 3'h0 : _GEN_571; // @[IoControl.scala 421:44 IoControl.scala 421:44]
  wire [2:0] _GEN_605 = 3'h1 == flush_head_idx ? 3'h0 : _GEN_572; // @[IoControl.scala 421:44 IoControl.scala 421:44]
  wire [2:0] _GEN_606 = 3'h2 == flush_head_idx ? 3'h0 : _GEN_573; // @[IoControl.scala 421:44 IoControl.scala 421:44]
  wire [2:0] _GEN_607 = 3'h3 == flush_head_idx ? 3'h0 : _GEN_574; // @[IoControl.scala 421:44 IoControl.scala 421:44]
  wire [2:0] _GEN_608 = 3'h4 == flush_head_idx ? 3'h0 : _GEN_575; // @[IoControl.scala 421:44 IoControl.scala 421:44]
  wire [2:0] _GEN_609 = 3'h5 == flush_head_idx ? 3'h0 : _GEN_576; // @[IoControl.scala 421:44 IoControl.scala 421:44]
  wire [2:0] _GEN_610 = 3'h6 == flush_head_idx ? 3'h0 : _GEN_577; // @[IoControl.scala 421:44 IoControl.scala 421:44]
  wire [2:0] _GEN_611 = 3'h7 == flush_head_idx ? 3'h0 : _GEN_578; // @[IoControl.scala 421:44 IoControl.scala 421:44]
  wire  _GEN_612 = 3'h0 == flush_head_idx ? 1'h0 : _GEN_579; // @[IoControl.scala 422:41 IoControl.scala 422:41]
  wire  _GEN_613 = 3'h1 == flush_head_idx ? 1'h0 : _GEN_580; // @[IoControl.scala 422:41 IoControl.scala 422:41]
  wire  _GEN_614 = 3'h2 == flush_head_idx ? 1'h0 : _GEN_581; // @[IoControl.scala 422:41 IoControl.scala 422:41]
  wire  _GEN_615 = 3'h3 == flush_head_idx ? 1'h0 : _GEN_582; // @[IoControl.scala 422:41 IoControl.scala 422:41]
  wire  _GEN_616 = 3'h4 == flush_head_idx ? 1'h0 : _GEN_583; // @[IoControl.scala 422:41 IoControl.scala 422:41]
  wire  _GEN_617 = 3'h5 == flush_head_idx ? 1'h0 : _GEN_584; // @[IoControl.scala 422:41 IoControl.scala 422:41]
  wire  _GEN_618 = 3'h6 == flush_head_idx ? 1'h0 : _GEN_585; // @[IoControl.scala 422:41 IoControl.scala 422:41]
  wire  _GEN_619 = 3'h7 == flush_head_idx ? 1'h0 : _GEN_586; // @[IoControl.scala 422:41 IoControl.scala 422:41]
  wire [2:0] _GEN_620 = _GEN_595 == io_rob_commit_0_bits_des_rob & io_rob_commit_0_valid & _GEN_603 ? _GEN_604 :
    _GEN_571; // @[IoControl.scala 420:138]
  wire [2:0] _GEN_621 = _GEN_595 == io_rob_commit_0_bits_des_rob & io_rob_commit_0_valid & _GEN_603 ? _GEN_605 :
    _GEN_572; // @[IoControl.scala 420:138]
  wire [2:0] _GEN_622 = _GEN_595 == io_rob_commit_0_bits_des_rob & io_rob_commit_0_valid & _GEN_603 ? _GEN_606 :
    _GEN_573; // @[IoControl.scala 420:138]
  wire [2:0] _GEN_623 = _GEN_595 == io_rob_commit_0_bits_des_rob & io_rob_commit_0_valid & _GEN_603 ? _GEN_607 :
    _GEN_574; // @[IoControl.scala 420:138]
  wire [2:0] _GEN_624 = _GEN_595 == io_rob_commit_0_bits_des_rob & io_rob_commit_0_valid & _GEN_603 ? _GEN_608 :
    _GEN_575; // @[IoControl.scala 420:138]
  wire [2:0] _GEN_625 = _GEN_595 == io_rob_commit_0_bits_des_rob & io_rob_commit_0_valid & _GEN_603 ? _GEN_609 :
    _GEN_576; // @[IoControl.scala 420:138]
  wire [2:0] _GEN_626 = _GEN_595 == io_rob_commit_0_bits_des_rob & io_rob_commit_0_valid & _GEN_603 ? _GEN_610 :
    _GEN_577; // @[IoControl.scala 420:138]
  wire [2:0] _GEN_627 = _GEN_595 == io_rob_commit_0_bits_des_rob & io_rob_commit_0_valid & _GEN_603 ? _GEN_611 :
    _GEN_578; // @[IoControl.scala 420:138]
  wire  _GEN_628 = _GEN_595 == io_rob_commit_0_bits_des_rob & io_rob_commit_0_valid & _GEN_603 ? _GEN_612 : _GEN_579; // @[IoControl.scala 420:138]
  wire  _GEN_629 = _GEN_595 == io_rob_commit_0_bits_des_rob & io_rob_commit_0_valid & _GEN_603 ? _GEN_613 : _GEN_580; // @[IoControl.scala 420:138]
  wire  _GEN_630 = _GEN_595 == io_rob_commit_0_bits_des_rob & io_rob_commit_0_valid & _GEN_603 ? _GEN_614 : _GEN_581; // @[IoControl.scala 420:138]
  wire  _GEN_631 = _GEN_595 == io_rob_commit_0_bits_des_rob & io_rob_commit_0_valid & _GEN_603 ? _GEN_615 : _GEN_582; // @[IoControl.scala 420:138]
  wire  _GEN_632 = _GEN_595 == io_rob_commit_0_bits_des_rob & io_rob_commit_0_valid & _GEN_603 ? _GEN_616 : _GEN_583; // @[IoControl.scala 420:138]
  wire  _GEN_633 = _GEN_595 == io_rob_commit_0_bits_des_rob & io_rob_commit_0_valid & _GEN_603 ? _GEN_617 : _GEN_584; // @[IoControl.scala 420:138]
  wire  _GEN_634 = _GEN_595 == io_rob_commit_0_bits_des_rob & io_rob_commit_0_valid & _GEN_603 ? _GEN_618 : _GEN_585; // @[IoControl.scala 420:138]
  wire  _GEN_635 = _GEN_595 == io_rob_commit_0_bits_des_rob & io_rob_commit_0_valid & _GEN_603 ? _GEN_619 : _GEN_586; // @[IoControl.scala 420:138]
  wire [2:0] _GEN_637 = 3'h0 == flush_head_idx ? 3'h0 : _GEN_620; // @[IoControl.scala 421:44 IoControl.scala 421:44]
  wire [2:0] _GEN_638 = 3'h1 == flush_head_idx ? 3'h0 : _GEN_621; // @[IoControl.scala 421:44 IoControl.scala 421:44]
  wire [2:0] _GEN_639 = 3'h2 == flush_head_idx ? 3'h0 : _GEN_622; // @[IoControl.scala 421:44 IoControl.scala 421:44]
  wire [2:0] _GEN_640 = 3'h3 == flush_head_idx ? 3'h0 : _GEN_623; // @[IoControl.scala 421:44 IoControl.scala 421:44]
  wire [2:0] _GEN_641 = 3'h4 == flush_head_idx ? 3'h0 : _GEN_624; // @[IoControl.scala 421:44 IoControl.scala 421:44]
  wire [2:0] _GEN_642 = 3'h5 == flush_head_idx ? 3'h0 : _GEN_625; // @[IoControl.scala 421:44 IoControl.scala 421:44]
  wire [2:0] _GEN_643 = 3'h6 == flush_head_idx ? 3'h0 : _GEN_626; // @[IoControl.scala 421:44 IoControl.scala 421:44]
  wire [2:0] _GEN_644 = 3'h7 == flush_head_idx ? 3'h0 : _GEN_627; // @[IoControl.scala 421:44 IoControl.scala 421:44]
  wire  _GEN_645 = 3'h0 == flush_head_idx ? 1'h0 : _GEN_628; // @[IoControl.scala 422:41 IoControl.scala 422:41]
  wire  _GEN_646 = 3'h1 == flush_head_idx ? 1'h0 : _GEN_629; // @[IoControl.scala 422:41 IoControl.scala 422:41]
  wire  _GEN_647 = 3'h2 == flush_head_idx ? 1'h0 : _GEN_630; // @[IoControl.scala 422:41 IoControl.scala 422:41]
  wire  _GEN_648 = 3'h3 == flush_head_idx ? 1'h0 : _GEN_631; // @[IoControl.scala 422:41 IoControl.scala 422:41]
  wire  _GEN_649 = 3'h4 == flush_head_idx ? 1'h0 : _GEN_632; // @[IoControl.scala 422:41 IoControl.scala 422:41]
  wire  _GEN_650 = 3'h5 == flush_head_idx ? 1'h0 : _GEN_633; // @[IoControl.scala 422:41 IoControl.scala 422:41]
  wire  _GEN_651 = 3'h6 == flush_head_idx ? 1'h0 : _GEN_634; // @[IoControl.scala 422:41 IoControl.scala 422:41]
  wire  _GEN_652 = 3'h7 == flush_head_idx ? 1'h0 : _GEN_635; // @[IoControl.scala 422:41 IoControl.scala 422:41]
  wire [2:0] _GEN_653 = _GEN_595 == io_rob_commit_1_bits_des_rob & io_rob_commit_1_valid & _GEN_603 ? _GEN_637 :
    _GEN_620; // @[IoControl.scala 420:138]
  wire [2:0] _GEN_654 = _GEN_595 == io_rob_commit_1_bits_des_rob & io_rob_commit_1_valid & _GEN_603 ? _GEN_638 :
    _GEN_621; // @[IoControl.scala 420:138]
  wire [2:0] _GEN_655 = _GEN_595 == io_rob_commit_1_bits_des_rob & io_rob_commit_1_valid & _GEN_603 ? _GEN_639 :
    _GEN_622; // @[IoControl.scala 420:138]
  wire [2:0] _GEN_656 = _GEN_595 == io_rob_commit_1_bits_des_rob & io_rob_commit_1_valid & _GEN_603 ? _GEN_640 :
    _GEN_623; // @[IoControl.scala 420:138]
  wire [2:0] _GEN_657 = _GEN_595 == io_rob_commit_1_bits_des_rob & io_rob_commit_1_valid & _GEN_603 ? _GEN_641 :
    _GEN_624; // @[IoControl.scala 420:138]
  wire [2:0] _GEN_658 = _GEN_595 == io_rob_commit_1_bits_des_rob & io_rob_commit_1_valid & _GEN_603 ? _GEN_642 :
    _GEN_625; // @[IoControl.scala 420:138]
  wire [2:0] _GEN_659 = _GEN_595 == io_rob_commit_1_bits_des_rob & io_rob_commit_1_valid & _GEN_603 ? _GEN_643 :
    _GEN_626; // @[IoControl.scala 420:138]
  wire [2:0] _GEN_660 = _GEN_595 == io_rob_commit_1_bits_des_rob & io_rob_commit_1_valid & _GEN_603 ? _GEN_644 :
    _GEN_627; // @[IoControl.scala 420:138]
  wire  _GEN_661 = _GEN_595 == io_rob_commit_1_bits_des_rob & io_rob_commit_1_valid & _GEN_603 ? _GEN_645 : _GEN_628; // @[IoControl.scala 420:138]
  wire  _GEN_662 = _GEN_595 == io_rob_commit_1_bits_des_rob & io_rob_commit_1_valid & _GEN_603 ? _GEN_646 : _GEN_629; // @[IoControl.scala 420:138]
  wire  _GEN_663 = _GEN_595 == io_rob_commit_1_bits_des_rob & io_rob_commit_1_valid & _GEN_603 ? _GEN_647 : _GEN_630; // @[IoControl.scala 420:138]
  wire  _GEN_664 = _GEN_595 == io_rob_commit_1_bits_des_rob & io_rob_commit_1_valid & _GEN_603 ? _GEN_648 : _GEN_631; // @[IoControl.scala 420:138]
  wire  _GEN_665 = _GEN_595 == io_rob_commit_1_bits_des_rob & io_rob_commit_1_valid & _GEN_603 ? _GEN_649 : _GEN_632; // @[IoControl.scala 420:138]
  wire  _GEN_666 = _GEN_595 == io_rob_commit_1_bits_des_rob & io_rob_commit_1_valid & _GEN_603 ? _GEN_650 : _GEN_633; // @[IoControl.scala 420:138]
  wire  _GEN_667 = _GEN_595 == io_rob_commit_1_bits_des_rob & io_rob_commit_1_valid & _GEN_603 ? _GEN_651 : _GEN_634; // @[IoControl.scala 420:138]
  wire  _GEN_668 = _GEN_595 == io_rob_commit_1_bits_des_rob & io_rob_commit_1_valid & _GEN_603 ? _GEN_652 : _GEN_635; // @[IoControl.scala 420:138]
  wire  will_drop_0 = _GEN_595 == io_rob_commit_1_bits_des_rob & io_rob_commit_1_valid & _GEN_603 | _GEN_595 ==
    io_rob_commit_0_bits_des_rob & io_rob_commit_0_valid & _GEN_603; // @[IoControl.scala 420:138 IoControl.scala 423:21]
  wire [6:0] flush_head_idx_hi_4 = uart_flush_head[6:0]; // @[IoControl.scala 106:12]
  wire  flush_head_idx_lo_4 = uart_flush_head[7]; // @[IoControl.scala 106:29]
  wire [7:0] _flush_head_idx_T_2 = {flush_head_idx_hi_4,flush_head_idx_lo_4}; // @[Cat.scala 30:58]
  wire [3:0] flush_head_idx_hi_5 = _flush_head_idx_T_2[7:4]; // @[OneHot.scala 30:18]
  wire [3:0] flush_head_idx_lo_5 = _flush_head_idx_T_2[3:0]; // @[OneHot.scala 31:18]
  wire  flush_head_idx_hi_6 = |flush_head_idx_hi_5; // @[OneHot.scala 32:14]
  wire [3:0] _flush_head_idx_T_3 = flush_head_idx_hi_5 | flush_head_idx_lo_5; // @[OneHot.scala 32:28]
  wire [1:0] flush_head_idx_hi_7 = _flush_head_idx_T_3[3:2]; // @[OneHot.scala 30:18]
  wire [1:0] flush_head_idx_lo_6 = _flush_head_idx_T_3[1:0]; // @[OneHot.scala 31:18]
  wire  flush_head_idx_hi_8 = |flush_head_idx_hi_7; // @[OneHot.scala 32:14]
  wire [1:0] _flush_head_idx_T_4 = flush_head_idx_hi_7 | flush_head_idx_lo_6; // @[OneHot.scala 32:28]
  wire  flush_head_idx_lo_7 = _flush_head_idx_T_4[1]; // @[CircuitMath.scala 30:8]
  wire [2:0] flush_head_idx_1 = {flush_head_idx_hi_6,flush_head_idx_hi_8,flush_head_idx_lo_7}; // @[Cat.scala 30:58]
  wire [2:0] _GEN_671 = 3'h1 == flush_head_idx_1 ? uart_buffer_1_rob_idx : uart_buffer_0_rob_idx; // @[IoControl.scala 420:47 IoControl.scala 420:47]
  wire [2:0] _GEN_672 = 3'h2 == flush_head_idx_1 ? uart_buffer_2_rob_idx : _GEN_671; // @[IoControl.scala 420:47 IoControl.scala 420:47]
  wire [2:0] _GEN_673 = 3'h3 == flush_head_idx_1 ? uart_buffer_3_rob_idx : _GEN_672; // @[IoControl.scala 420:47 IoControl.scala 420:47]
  wire [2:0] _GEN_674 = 3'h4 == flush_head_idx_1 ? uart_buffer_4_rob_idx : _GEN_673; // @[IoControl.scala 420:47 IoControl.scala 420:47]
  wire [2:0] _GEN_675 = 3'h5 == flush_head_idx_1 ? uart_buffer_5_rob_idx : _GEN_674; // @[IoControl.scala 420:47 IoControl.scala 420:47]
  wire [2:0] _GEN_676 = 3'h6 == flush_head_idx_1 ? uart_buffer_6_rob_idx : _GEN_675; // @[IoControl.scala 420:47 IoControl.scala 420:47]
  wire [2:0] _GEN_677 = 3'h7 == flush_head_idx_1 ? uart_buffer_7_rob_idx : _GEN_676; // @[IoControl.scala 420:47 IoControl.scala 420:47]
  wire  _GEN_679 = 3'h1 == flush_head_idx_1 ? uart_buffer_wait_1 : uart_buffer_wait_0; // @[IoControl.scala 420:103 IoControl.scala 420:103]
  wire  _GEN_680 = 3'h2 == flush_head_idx_1 ? uart_buffer_wait_2 : _GEN_679; // @[IoControl.scala 420:103 IoControl.scala 420:103]
  wire  _GEN_681 = 3'h3 == flush_head_idx_1 ? uart_buffer_wait_3 : _GEN_680; // @[IoControl.scala 420:103 IoControl.scala 420:103]
  wire  _GEN_682 = 3'h4 == flush_head_idx_1 ? uart_buffer_wait_4 : _GEN_681; // @[IoControl.scala 420:103 IoControl.scala 420:103]
  wire  _GEN_683 = 3'h5 == flush_head_idx_1 ? uart_buffer_wait_5 : _GEN_682; // @[IoControl.scala 420:103 IoControl.scala 420:103]
  wire  _GEN_684 = 3'h6 == flush_head_idx_1 ? uart_buffer_wait_6 : _GEN_683; // @[IoControl.scala 420:103 IoControl.scala 420:103]
  wire  _GEN_685 = 3'h7 == flush_head_idx_1 ? uart_buffer_wait_7 : _GEN_684; // @[IoControl.scala 420:103 IoControl.scala 420:103]
  wire [2:0] _GEN_686 = 3'h0 == flush_head_idx_1 ? 3'h0 : _GEN_653; // @[IoControl.scala 421:44 IoControl.scala 421:44]
  wire [2:0] _GEN_687 = 3'h1 == flush_head_idx_1 ? 3'h0 : _GEN_654; // @[IoControl.scala 421:44 IoControl.scala 421:44]
  wire [2:0] _GEN_688 = 3'h2 == flush_head_idx_1 ? 3'h0 : _GEN_655; // @[IoControl.scala 421:44 IoControl.scala 421:44]
  wire [2:0] _GEN_689 = 3'h3 == flush_head_idx_1 ? 3'h0 : _GEN_656; // @[IoControl.scala 421:44 IoControl.scala 421:44]
  wire [2:0] _GEN_690 = 3'h4 == flush_head_idx_1 ? 3'h0 : _GEN_657; // @[IoControl.scala 421:44 IoControl.scala 421:44]
  wire [2:0] _GEN_691 = 3'h5 == flush_head_idx_1 ? 3'h0 : _GEN_658; // @[IoControl.scala 421:44 IoControl.scala 421:44]
  wire [2:0] _GEN_692 = 3'h6 == flush_head_idx_1 ? 3'h0 : _GEN_659; // @[IoControl.scala 421:44 IoControl.scala 421:44]
  wire [2:0] _GEN_693 = 3'h7 == flush_head_idx_1 ? 3'h0 : _GEN_660; // @[IoControl.scala 421:44 IoControl.scala 421:44]
  wire  _GEN_694 = 3'h0 == flush_head_idx_1 ? 1'h0 : _GEN_661; // @[IoControl.scala 422:41 IoControl.scala 422:41]
  wire  _GEN_695 = 3'h1 == flush_head_idx_1 ? 1'h0 : _GEN_662; // @[IoControl.scala 422:41 IoControl.scala 422:41]
  wire  _GEN_696 = 3'h2 == flush_head_idx_1 ? 1'h0 : _GEN_663; // @[IoControl.scala 422:41 IoControl.scala 422:41]
  wire  _GEN_697 = 3'h3 == flush_head_idx_1 ? 1'h0 : _GEN_664; // @[IoControl.scala 422:41 IoControl.scala 422:41]
  wire  _GEN_698 = 3'h4 == flush_head_idx_1 ? 1'h0 : _GEN_665; // @[IoControl.scala 422:41 IoControl.scala 422:41]
  wire  _GEN_699 = 3'h5 == flush_head_idx_1 ? 1'h0 : _GEN_666; // @[IoControl.scala 422:41 IoControl.scala 422:41]
  wire  _GEN_700 = 3'h6 == flush_head_idx_1 ? 1'h0 : _GEN_667; // @[IoControl.scala 422:41 IoControl.scala 422:41]
  wire  _GEN_701 = 3'h7 == flush_head_idx_1 ? 1'h0 : _GEN_668; // @[IoControl.scala 422:41 IoControl.scala 422:41]
  wire [2:0] _GEN_702 = _GEN_677 == io_rob_commit_0_bits_des_rob & io_rob_commit_0_valid & _GEN_685 ? _GEN_686 :
    _GEN_653; // @[IoControl.scala 420:138]
  wire [2:0] _GEN_703 = _GEN_677 == io_rob_commit_0_bits_des_rob & io_rob_commit_0_valid & _GEN_685 ? _GEN_687 :
    _GEN_654; // @[IoControl.scala 420:138]
  wire [2:0] _GEN_704 = _GEN_677 == io_rob_commit_0_bits_des_rob & io_rob_commit_0_valid & _GEN_685 ? _GEN_688 :
    _GEN_655; // @[IoControl.scala 420:138]
  wire [2:0] _GEN_705 = _GEN_677 == io_rob_commit_0_bits_des_rob & io_rob_commit_0_valid & _GEN_685 ? _GEN_689 :
    _GEN_656; // @[IoControl.scala 420:138]
  wire [2:0] _GEN_706 = _GEN_677 == io_rob_commit_0_bits_des_rob & io_rob_commit_0_valid & _GEN_685 ? _GEN_690 :
    _GEN_657; // @[IoControl.scala 420:138]
  wire [2:0] _GEN_707 = _GEN_677 == io_rob_commit_0_bits_des_rob & io_rob_commit_0_valid & _GEN_685 ? _GEN_691 :
    _GEN_658; // @[IoControl.scala 420:138]
  wire [2:0] _GEN_708 = _GEN_677 == io_rob_commit_0_bits_des_rob & io_rob_commit_0_valid & _GEN_685 ? _GEN_692 :
    _GEN_659; // @[IoControl.scala 420:138]
  wire [2:0] _GEN_709 = _GEN_677 == io_rob_commit_0_bits_des_rob & io_rob_commit_0_valid & _GEN_685 ? _GEN_693 :
    _GEN_660; // @[IoControl.scala 420:138]
  wire  _GEN_710 = _GEN_677 == io_rob_commit_0_bits_des_rob & io_rob_commit_0_valid & _GEN_685 ? _GEN_694 : _GEN_661; // @[IoControl.scala 420:138]
  wire  _GEN_711 = _GEN_677 == io_rob_commit_0_bits_des_rob & io_rob_commit_0_valid & _GEN_685 ? _GEN_695 : _GEN_662; // @[IoControl.scala 420:138]
  wire  _GEN_712 = _GEN_677 == io_rob_commit_0_bits_des_rob & io_rob_commit_0_valid & _GEN_685 ? _GEN_696 : _GEN_663; // @[IoControl.scala 420:138]
  wire  _GEN_713 = _GEN_677 == io_rob_commit_0_bits_des_rob & io_rob_commit_0_valid & _GEN_685 ? _GEN_697 : _GEN_664; // @[IoControl.scala 420:138]
  wire  _GEN_714 = _GEN_677 == io_rob_commit_0_bits_des_rob & io_rob_commit_0_valid & _GEN_685 ? _GEN_698 : _GEN_665; // @[IoControl.scala 420:138]
  wire  _GEN_715 = _GEN_677 == io_rob_commit_0_bits_des_rob & io_rob_commit_0_valid & _GEN_685 ? _GEN_699 : _GEN_666; // @[IoControl.scala 420:138]
  wire  _GEN_716 = _GEN_677 == io_rob_commit_0_bits_des_rob & io_rob_commit_0_valid & _GEN_685 ? _GEN_700 : _GEN_667; // @[IoControl.scala 420:138]
  wire  _GEN_717 = _GEN_677 == io_rob_commit_0_bits_des_rob & io_rob_commit_0_valid & _GEN_685 ? _GEN_701 : _GEN_668; // @[IoControl.scala 420:138]
  wire  will_drop_1 = _GEN_677 == io_rob_commit_1_bits_des_rob & io_rob_commit_1_valid & _GEN_685 | _GEN_677 ==
    io_rob_commit_0_bits_des_rob & io_rob_commit_0_valid & _GEN_685; // @[IoControl.scala 420:138 IoControl.scala 423:21]
  wire [5:0] next_flush_head_hi_1 = uart_flush_head[5:0]; // @[IoControl.scala 106:12]
  wire [1:0] next_flush_head_lo_1 = uart_flush_head[7:6]; // @[IoControl.scala 106:29]
  wire [7:0] _next_flush_head_T_2 = {next_flush_head_hi_1,next_flush_head_lo_1}; // @[Cat.scala 30:58]
  wire  _GEN_752 = will_drop_0 | will_drop_1 ? 1'h0 : maybe_true_full; // @[IoControl.scala 432:36 IoControl.scala 433:20 IoControl.scala 386:32]
  wire  _GEN_753 = uart_enq | _GEN_752; // @[IoControl.scala 430:17 IoControl.scala 431:20]
  wire  _GEN_754 = uart_deq ? 1'h0 : maybe_full; // @[IoControl.scala 437:23 IoControl.scala 438:15 IoControl.scala 385:27]
  wire  _GEN_755 = uart_enq | _GEN_754; // @[IoControl.scala 435:17 IoControl.scala 436:15]
  reg  txd_uart_start; // @[IoControl.scala 453:31]
  reg [7:0] txd_uart_data; // @[IoControl.scala 454:30]
  wire [31:0] _dcache_buffer_T = {24'h0,read_data}; // @[Cat.scala 30:58]
  wire [31:0] _dcache_buffer_T_1 = {30'h0,_uart_deq_T,_T_57}; // @[Cat.scala 30:58]
  wire [31:0] _GEN_768 = dcache_read_uart_state ? _dcache_buffer_T_1 : _GEN_511; // @[IoControl.scala 481:41 IoControl.scala 482:22]
  wire  _GEN_769 = dcache_read_uart_state | _GEN_512; // @[IoControl.scala 481:41 IoControl.scala 483:26]
  wire [1:0] _GEN_770 = dcache_read_uart_state ? 2'h1 : uart_state; // @[IoControl.scala 481:41 IoControl.scala 484:19 IoControl.scala 452:27]
  wire  _GEN_772 = dcache_read_uart & _uart_deq_T | _GEN_769; // @[IoControl.scala 475:48 IoControl.scala 477:26]
  wire  _GEN_776 = dcache_write_uart & ~io_txd_uart_busy | txd_uart_start; // @[IoControl.scala 470:50 IoControl.scala 471:23 IoControl.scala 453:31]
  wire  _GEN_778 = dcache_write_uart & ~io_txd_uart_busy | _GEN_513; // @[IoControl.scala 470:50 IoControl.scala 473:30]
  wire  _T_60 = 2'h2 == uart_state; // @[Conditional.scala 37:30]
  wire  _T_61 = 2'h1 == uart_state; // @[Conditional.scala 37:30]
  assign io_icache_read_req_ready = icache_data_valid; // @[IoControl.scala 157:28]
  assign io_icache_read_resp_bits_data = {io_icache_read_resp_bits_data_hi,io_icache_read_resp_bits_data_lo}; // @[IoControl.scala 159:56]
  assign io_dcache_read_req_ready = dcache_data_valid; // @[IoControl.scala 162:28]
  assign io_dcache_read_resp_bits_data = dcache_buffer; // @[IoControl.scala 164:33]
  assign io_dcache_write_req_ready = _T_56 ? _GEN_778 : _GEN_513; // @[Conditional.scala 40:58]
  assign io_base_ram_ctrl_ctrl_data_out = base_ram_ctrl_data_out; // @[IoControl.scala 116:25]
  assign io_base_ram_ctrl_ctrl_addr = base_ram_ctrl_addr; // @[IoControl.scala 116:25]
  assign io_base_ram_ctrl_ctrl_be_n = base_ram_ctrl_be_n; // @[IoControl.scala 116:25]
  assign io_base_ram_ctrl_ctrl_ce_n = base_ram_ctrl_ce_n; // @[IoControl.scala 116:25]
  assign io_base_ram_ctrl_ctrl_oe_n = base_ram_ctrl_oe_n; // @[IoControl.scala 116:25]
  assign io_base_ram_ctrl_ctrl_we_n = base_ram_ctrl_we_n; // @[IoControl.scala 116:25]
  assign io_ext_ram_ctrl_ctrl_data_out = ext_ram_ctrl_data_out; // @[IoControl.scala 117:24]
  assign io_ext_ram_ctrl_ctrl_addr = ext_ram_ctrl_addr; // @[IoControl.scala 117:24]
  assign io_ext_ram_ctrl_ctrl_be_n = ext_ram_ctrl_be_n; // @[IoControl.scala 117:24]
  assign io_ext_ram_ctrl_ctrl_ce_n = ext_ram_ctrl_ce_n; // @[IoControl.scala 117:24]
  assign io_ext_ram_ctrl_ctrl_oe_n = ext_ram_ctrl_oe_n; // @[IoControl.scala 117:24]
  assign io_ext_ram_ctrl_ctrl_we_n = ext_ram_ctrl_we_n; // @[IoControl.scala 117:24]
  assign io_rxd_uart_clear = io_rxd_uart_ready & _uart_enq_T; // @[IoControl.scala 458:25]
  assign io_txd_uart_start = txd_uart_start; // @[IoControl.scala 455:20]
  assign io_txd_uart_data = txd_uart_data; // @[IoControl.scala 456:19]
  assign io_debug_base_state = base_state; // @[IoControl.scala 143:23]
  assign io_debug_icache_read_base = io_icache_read_req_bits_addr[31:22] == 10'h200 & io_icache_read_req_valid; // @[IoControl.scala 127:101]
  assign io_debug_icache_read_ext = io_icache_read_req_bits_addr[31:22] == 10'h201 & io_icache_read_req_valid; // @[IoControl.scala 128:101]
  assign io_debug_dcache_read_base = io_dcache_read_req_bits_addr[31:22] == 10'h200 & io_dcache_read_req_valid; // @[IoControl.scala 129:101]
  assign io_debug_dcache_read_ext = io_dcache_read_req_bits_addr[31:22] == 10'h201 & io_dcache_read_req_valid; // @[IoControl.scala 130:101]
  assign io_debug_dcache_write_base = io_dcache_write_req_bits_addr[31:22] == 10'h200 & io_dcache_write_req_valid; // @[IoControl.scala 131:102]
  assign io_debug_dcache_write_ext = io_dcache_write_req_bits_addr[31:22] == 10'h201 & io_dcache_write_req_valid; // @[IoControl.scala 132:102]
  assign io_debug_icache_read_addr = io_icache_read_req_bits_addr[21:2]; // @[IoControl.scala 136:67]
  assign io_debug_dcache_read_addr = io_dcache_read_req_bits_addr[21:2]; // @[IoControl.scala 137:67]
  assign io_debug_dcache_write_addr = io_dcache_write_req_bits_addr[21:2]; // @[IoControl.scala 138:68]
  always @(posedge clock) begin
    if (reset) begin // @[IoControl.scala 498:24]
      base_ram_ctrl_data_out <= 32'h0; // @[IoControl.scala 12:14]
    end else if (_T_4) begin // @[Conditional.scala 40:58]
      if (dcache_write_base) begin // @[IoControl.scala 206:31]
        base_ram_ctrl_data_out <= io_dcache_write_req_bits_data; // @[IoControl.scala 30:14]
      end else if (dcache_read_base) begin // @[IoControl.scala 212:36]
        base_ram_ctrl_data_out <= 32'h0; // @[IoControl.scala 21:14]
      end else begin
        base_ram_ctrl_data_out <= _GEN_35;
      end
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      if (_icache_read_other_T) begin // @[IoControl.scala 225:31]
        base_ram_ctrl_data_out <= 32'h0; // @[IoControl.scala 12:14]
      end else begin
        base_ram_ctrl_data_out <= _GEN_118;
      end
    end else if (!(_T_15)) begin // @[Conditional.scala 39:67]
      base_ram_ctrl_data_out <= _GEN_207;
    end
    if (reset) begin // @[IoControl.scala 498:24]
      base_ram_ctrl_addr <= 20'h0; // @[IoControl.scala 13:10]
    end else if (_T_4) begin // @[Conditional.scala 40:58]
      if (dcache_write_base) begin // @[IoControl.scala 206:31]
        base_ram_ctrl_addr <= dcache_write_addr; // @[IoControl.scala 31:10]
      end else if (dcache_read_base) begin // @[IoControl.scala 212:36]
        base_ram_ctrl_addr <= dcache_read_addr; // @[IoControl.scala 22:10]
      end else begin
        base_ram_ctrl_addr <= _GEN_36;
      end
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      if (_icache_read_other_T) begin // @[IoControl.scala 225:31]
        base_ram_ctrl_addr <= 20'h0; // @[IoControl.scala 13:10]
      end else begin
        base_ram_ctrl_addr <= _GEN_119;
      end
    end else if (!(_T_15)) begin // @[Conditional.scala 39:67]
      base_ram_ctrl_addr <= _GEN_208;
    end
    if (reset) begin // @[IoControl.scala 498:24]
      base_ram_ctrl_be_n <= 4'hf; // @[IoControl.scala 14:10]
    end else if (_T_4) begin // @[Conditional.scala 40:58]
      if (dcache_write_base) begin // @[IoControl.scala 206:31]
        base_ram_ctrl_be_n <= _T_5; // @[IoControl.scala 32:10]
      end else if (dcache_read_base) begin // @[IoControl.scala 212:36]
        base_ram_ctrl_be_n <= 4'h0; // @[IoControl.scala 23:10]
      end else begin
        base_ram_ctrl_be_n <= _GEN_37;
      end
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      if (_icache_read_other_T) begin // @[IoControl.scala 225:31]
        base_ram_ctrl_be_n <= 4'hf; // @[IoControl.scala 14:10]
      end else begin
        base_ram_ctrl_be_n <= _GEN_120;
      end
    end else if (!(_T_15)) begin // @[Conditional.scala 39:67]
      base_ram_ctrl_be_n <= _GEN_209;
    end
    base_ram_ctrl_ce_n <= reset | _GEN_257; // @[IoControl.scala 498:24 IoControl.scala 15:10]
    base_ram_ctrl_oe_n <= reset | _GEN_258; // @[IoControl.scala 498:24 IoControl.scala 16:10]
    base_ram_ctrl_we_n <= reset | _GEN_259; // @[IoControl.scala 498:24 IoControl.scala 17:10]
    if (reset) begin // @[IoControl.scala 498:24]
      ext_ram_ctrl_data_out <= 32'h0; // @[IoControl.scala 12:14]
    end else if (_T_23) begin // @[Conditional.scala 40:58]
      if (dcache_read_ext) begin // @[IoControl.scala 292:29]
        ext_ram_ctrl_data_out <= 32'h0; // @[IoControl.scala 21:14]
      end else if (dcache_write_ext) begin // @[IoControl.scala 297:36]
        ext_ram_ctrl_data_out <= io_dcache_write_req_bits_data; // @[IoControl.scala 30:14]
      end else begin
        ext_ram_ctrl_data_out <= _GEN_275;
      end
    end else if (_T_25) begin // @[Conditional.scala 39:67]
      if (_icache_read_other_T_1) begin // @[IoControl.scala 311:30]
        ext_ram_ctrl_data_out <= 32'h0; // @[IoControl.scala 12:14]
      end else begin
        ext_ram_ctrl_data_out <= _GEN_358;
      end
    end else if (!(_T_34)) begin // @[Conditional.scala 39:67]
      ext_ram_ctrl_data_out <= _GEN_447;
    end
    if (reset) begin // @[IoControl.scala 498:24]
      ext_ram_ctrl_addr <= 20'h0; // @[IoControl.scala 13:10]
    end else if (_T_23) begin // @[Conditional.scala 40:58]
      if (dcache_read_ext) begin // @[IoControl.scala 292:29]
        ext_ram_ctrl_addr <= dcache_read_addr; // @[IoControl.scala 22:10]
      end else if (dcache_write_ext) begin // @[IoControl.scala 297:36]
        ext_ram_ctrl_addr <= dcache_write_addr; // @[IoControl.scala 31:10]
      end else begin
        ext_ram_ctrl_addr <= _GEN_276;
      end
    end else if (_T_25) begin // @[Conditional.scala 39:67]
      if (_icache_read_other_T_1) begin // @[IoControl.scala 311:30]
        ext_ram_ctrl_addr <= 20'h0; // @[IoControl.scala 13:10]
      end else begin
        ext_ram_ctrl_addr <= _GEN_359;
      end
    end else if (!(_T_34)) begin // @[Conditional.scala 39:67]
      ext_ram_ctrl_addr <= _GEN_448;
    end
    if (reset) begin // @[IoControl.scala 498:24]
      ext_ram_ctrl_be_n <= 4'hf; // @[IoControl.scala 14:10]
    end else if (_T_23) begin // @[Conditional.scala 40:58]
      if (dcache_read_ext) begin // @[IoControl.scala 292:29]
        ext_ram_ctrl_be_n <= 4'h0; // @[IoControl.scala 23:10]
      end else if (dcache_write_ext) begin // @[IoControl.scala 297:36]
        ext_ram_ctrl_be_n <= _T_5; // @[IoControl.scala 32:10]
      end else begin
        ext_ram_ctrl_be_n <= _GEN_277;
      end
    end else if (_T_25) begin // @[Conditional.scala 39:67]
      if (_icache_read_other_T_1) begin // @[IoControl.scala 311:30]
        ext_ram_ctrl_be_n <= 4'hf; // @[IoControl.scala 14:10]
      end else begin
        ext_ram_ctrl_be_n <= _GEN_360;
      end
    end else if (!(_T_34)) begin // @[Conditional.scala 39:67]
      ext_ram_ctrl_be_n <= _GEN_449;
    end
    ext_ram_ctrl_ce_n <= reset | _GEN_497; // @[IoControl.scala 498:24 IoControl.scala 15:10]
    ext_ram_ctrl_oe_n <= reset | _GEN_498; // @[IoControl.scala 498:24 IoControl.scala 16:10]
    ext_ram_ctrl_we_n <= reset | _GEN_499; // @[IoControl.scala 498:24 IoControl.scala 17:10]
    if (reset) begin // @[IoControl.scala 120:46]
      base_state <= 3'h0; // @[IoControl.scala 120:46]
    end else if (_T_4) begin // @[Conditional.scala 40:58]
      if (dcache_write_base) begin // @[IoControl.scala 206:31]
        base_state <= 3'h3; // @[IoControl.scala 207:20]
      end else if (dcache_read_base) begin // @[IoControl.scala 212:36]
        base_state <= 3'h2; // @[IoControl.scala 213:20]
      end else begin
        base_state <= _GEN_34;
      end
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      if (_icache_read_other_T) begin // @[IoControl.scala 225:31]
        base_state <= 3'h0; // @[IoControl.scala 227:20]
      end else begin
        base_state <= _GEN_125;
      end
    end else if (_T_15) begin // @[Conditional.scala 39:67]
      base_state <= 3'h0; // @[IoControl.scala 252:20]
    end else begin
      base_state <= _GEN_213;
    end
    if (reset) begin // @[IoControl.scala 121:46]
      base_clock_counter <= 4'h0; // @[IoControl.scala 121:46]
    end else if (_T_4) begin // @[Conditional.scala 40:58]
      if (dcache_write_base) begin // @[IoControl.scala 206:31]
        base_clock_counter <= 4'h0; // @[IoControl.scala 210:28]
      end else if (dcache_read_base) begin // @[IoControl.scala 212:36]
        base_clock_counter <= 4'h0; // @[IoControl.scala 215:28]
      end else begin
        base_clock_counter <= _GEN_41;
      end
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      if (_icache_read_other_T) begin // @[IoControl.scala 225:31]
        base_clock_counter <= 4'h0; // @[IoControl.scala 228:28]
      end else begin
        base_clock_counter <= _GEN_127;
      end
    end else if (!(_T_15)) begin // @[Conditional.scala 39:67]
      base_clock_counter <= _GEN_214;
    end
    if (reset) begin // @[IoControl.scala 122:45]
      base_wait_counter <= 4'h0; // @[IoControl.scala 122:45]
    end else if (_T_4) begin // @[Conditional.scala 40:58]
      if (dcache_write_base) begin // @[IoControl.scala 206:31]
        base_wait_counter <= 4'h0; // @[IoControl.scala 211:27]
      end else if (dcache_read_base) begin // @[IoControl.scala 212:36]
        base_wait_counter <= 4'h0; // @[IoControl.scala 216:27]
      end else begin
        base_wait_counter <= _GEN_42;
      end
    end else if (_T_6) begin // @[Conditional.scala 39:67]
      if (_icache_read_other_T) begin // @[IoControl.scala 225:31]
        base_wait_counter <= 4'h0; // @[IoControl.scala 229:27]
      end else begin
        base_wait_counter <= _GEN_126;
      end
    end else if (!(_T_15)) begin // @[Conditional.scala 39:67]
      base_wait_counter <= _GEN_215;
    end
    if (reset) begin // @[IoControl.scala 123:46]
      ext_state <= 3'h0; // @[IoControl.scala 123:46]
    end else if (_T_23) begin // @[Conditional.scala 40:58]
      if (dcache_read_ext) begin // @[IoControl.scala 292:29]
        ext_state <= 3'h2; // @[IoControl.scala 293:19]
      end else if (dcache_write_ext) begin // @[IoControl.scala 297:36]
        ext_state <= 3'h3; // @[IoControl.scala 298:19]
      end else begin
        ext_state <= _GEN_274;
      end
    end else if (_T_25) begin // @[Conditional.scala 39:67]
      if (_icache_read_other_T_1) begin // @[IoControl.scala 311:30]
        ext_state <= 3'h0; // @[IoControl.scala 313:19]
      end else begin
        ext_state <= _GEN_365;
      end
    end else if (_T_34) begin // @[Conditional.scala 39:67]
      ext_state <= 3'h0; // @[IoControl.scala 338:17]
    end else begin
      ext_state <= _GEN_453;
    end
    if (reset) begin // @[IoControl.scala 124:46]
      ext_clock_counter <= 4'h0; // @[IoControl.scala 124:46]
    end else if (_T_23) begin // @[Conditional.scala 40:58]
      if (dcache_read_ext) begin // @[IoControl.scala 292:29]
        ext_clock_counter <= 4'h0; // @[IoControl.scala 295:27]
      end else if (dcache_write_ext) begin // @[IoControl.scala 297:36]
        ext_clock_counter <= 4'h0; // @[IoControl.scala 301:27]
      end else begin
        ext_clock_counter <= _GEN_281;
      end
    end else if (_T_25) begin // @[Conditional.scala 39:67]
      if (_icache_read_other_T_1) begin // @[IoControl.scala 311:30]
        ext_clock_counter <= 4'h0; // @[IoControl.scala 314:27]
      end else begin
        ext_clock_counter <= _GEN_367;
      end
    end else if (!(_T_34)) begin // @[Conditional.scala 39:67]
      ext_clock_counter <= _GEN_454;
    end
    if (reset) begin // @[IoControl.scala 125:45]
      ext_wait_counter <= 4'h0; // @[IoControl.scala 125:45]
    end else if (_T_23) begin // @[Conditional.scala 40:58]
      if (dcache_read_ext) begin // @[IoControl.scala 292:29]
        ext_wait_counter <= 4'h0; // @[IoControl.scala 296:26]
      end else if (dcache_write_ext) begin // @[IoControl.scala 297:36]
        ext_wait_counter <= 4'h0; // @[IoControl.scala 302:26]
      end else begin
        ext_wait_counter <= _GEN_282;
      end
    end else if (_T_25) begin // @[Conditional.scala 39:67]
      if (_icache_read_other_T_1) begin // @[IoControl.scala 311:30]
        ext_wait_counter <= 4'h0; // @[IoControl.scala 315:26]
      end else begin
        ext_wait_counter <= _GEN_366;
      end
    end else if (!(_T_34)) begin // @[Conditional.scala 39:67]
      ext_wait_counter <= _GEN_455;
    end
    if (reset) begin // @[IoControl.scala 155:34]
      icache_buffer_0 <= 32'h0; // @[IoControl.scala 155:34]
    end else if (_T_23) begin // @[Conditional.scala 40:58]
      icache_buffer_0 <= _GEN_262;
    end else if (_T_25) begin // @[Conditional.scala 39:67]
      if (_icache_read_other_T_1) begin // @[IoControl.scala 311:30]
        icache_buffer_0 <= _GEN_262;
      end else begin
        icache_buffer_0 <= _GEN_350;
      end
    end else begin
      icache_buffer_0 <= _GEN_262;
    end
    if (reset) begin // @[IoControl.scala 155:34]
      icache_buffer_1 <= 32'h0; // @[IoControl.scala 155:34]
    end else if (_T_23) begin // @[Conditional.scala 40:58]
      icache_buffer_1 <= _GEN_263;
    end else if (_T_25) begin // @[Conditional.scala 39:67]
      if (_icache_read_other_T_1) begin // @[IoControl.scala 311:30]
        icache_buffer_1 <= _GEN_263;
      end else begin
        icache_buffer_1 <= _GEN_351;
      end
    end else begin
      icache_buffer_1 <= _GEN_263;
    end
    if (reset) begin // @[IoControl.scala 155:34]
      icache_buffer_2 <= 32'h0; // @[IoControl.scala 155:34]
    end else if (_T_23) begin // @[Conditional.scala 40:58]
      icache_buffer_2 <= _GEN_264;
    end else if (_T_25) begin // @[Conditional.scala 39:67]
      if (_icache_read_other_T_1) begin // @[IoControl.scala 311:30]
        icache_buffer_2 <= _GEN_264;
      end else begin
        icache_buffer_2 <= _GEN_352;
      end
    end else begin
      icache_buffer_2 <= _GEN_264;
    end
    if (reset) begin // @[IoControl.scala 155:34]
      icache_buffer_3 <= 32'h0; // @[IoControl.scala 155:34]
    end else if (_T_23) begin // @[Conditional.scala 40:58]
      icache_buffer_3 <= _GEN_265;
    end else if (_T_25) begin // @[Conditional.scala 39:67]
      if (_icache_read_other_T_1) begin // @[IoControl.scala 311:30]
        icache_buffer_3 <= _GEN_265;
      end else begin
        icache_buffer_3 <= _GEN_353;
      end
    end else begin
      icache_buffer_3 <= _GEN_265;
    end
    if (reset) begin // @[IoControl.scala 155:34]
      icache_buffer_4 <= 32'h0; // @[IoControl.scala 155:34]
    end else if (_T_23) begin // @[Conditional.scala 40:58]
      icache_buffer_4 <= _GEN_266;
    end else if (_T_25) begin // @[Conditional.scala 39:67]
      if (_icache_read_other_T_1) begin // @[IoControl.scala 311:30]
        icache_buffer_4 <= _GEN_266;
      end else begin
        icache_buffer_4 <= _GEN_354;
      end
    end else begin
      icache_buffer_4 <= _GEN_266;
    end
    if (reset) begin // @[IoControl.scala 155:34]
      icache_buffer_5 <= 32'h0; // @[IoControl.scala 155:34]
    end else if (_T_23) begin // @[Conditional.scala 40:58]
      icache_buffer_5 <= _GEN_267;
    end else if (_T_25) begin // @[Conditional.scala 39:67]
      if (_icache_read_other_T_1) begin // @[IoControl.scala 311:30]
        icache_buffer_5 <= _GEN_267;
      end else begin
        icache_buffer_5 <= _GEN_355;
      end
    end else begin
      icache_buffer_5 <= _GEN_267;
    end
    if (reset) begin // @[IoControl.scala 155:34]
      icache_buffer_6 <= 32'h0; // @[IoControl.scala 155:34]
    end else if (_T_23) begin // @[Conditional.scala 40:58]
      icache_buffer_6 <= _GEN_268;
    end else if (_T_25) begin // @[Conditional.scala 39:67]
      if (_icache_read_other_T_1) begin // @[IoControl.scala 311:30]
        icache_buffer_6 <= _GEN_268;
      end else begin
        icache_buffer_6 <= _GEN_356;
      end
    end else begin
      icache_buffer_6 <= _GEN_268;
    end
    if (reset) begin // @[IoControl.scala 155:34]
      icache_buffer_7 <= 32'h0; // @[IoControl.scala 155:34]
    end else if (_T_23) begin // @[Conditional.scala 40:58]
      icache_buffer_7 <= _GEN_269;
    end else if (_T_25) begin // @[Conditional.scala 39:67]
      if (_icache_read_other_T_1) begin // @[IoControl.scala 311:30]
        icache_buffer_7 <= _GEN_269;
      end else begin
        icache_buffer_7 <= _GEN_357;
      end
    end else begin
      icache_buffer_7 <= _GEN_269;
    end
    if (reset) begin // @[IoControl.scala 156:34]
      icache_data_valid <= 1'h0; // @[IoControl.scala 156:34]
    end else if (_T_23) begin // @[Conditional.scala 40:58]
      icache_data_valid <= _GEN_270;
    end else if (_T_25) begin // @[Conditional.scala 39:67]
      if (_icache_read_other_T_1) begin // @[IoControl.scala 311:30]
        icache_data_valid <= _GEN_270;
      end else begin
        icache_data_valid <= _GEN_364;
      end
    end else if (_T_34) begin // @[Conditional.scala 39:67]
      icache_data_valid <= 1'h0; // @[IoControl.scala 339:25]
    end else begin
      icache_data_valid <= _GEN_270;
    end
    if (reset) begin // @[IoControl.scala 160:34]
      dcache_buffer <= 32'h0; // @[IoControl.scala 160:34]
    end else if (_T_56) begin // @[Conditional.scala 40:58]
      if (dcache_write_uart & ~io_txd_uart_busy) begin // @[IoControl.scala 470:50]
        dcache_buffer <= _GEN_511;
      end else if (dcache_read_uart & _uart_deq_T) begin // @[IoControl.scala 475:48]
        dcache_buffer <= _dcache_buffer_T; // @[IoControl.scala 476:22]
      end else begin
        dcache_buffer <= _GEN_768;
      end
    end else begin
      dcache_buffer <= _GEN_511;
    end
    if (reset) begin // @[IoControl.scala 161:34]
      dcache_data_valid <= 1'h0; // @[IoControl.scala 161:34]
    end else if (_T_56) begin // @[Conditional.scala 40:58]
      if (dcache_write_uart & ~io_txd_uart_busy) begin // @[IoControl.scala 470:50]
        dcache_data_valid <= _GEN_512;
      end else begin
        dcache_data_valid <= _GEN_772;
      end
    end else if (_T_60) begin // @[Conditional.scala 39:67]
      dcache_data_valid <= _GEN_512;
    end else if (_T_61) begin // @[Conditional.scala 39:67]
      dcache_data_valid <= 1'h0; // @[IoControl.scala 492:24]
    end else begin
      dcache_data_valid <= _GEN_512;
    end
    if (reset) begin // @[IoControl.scala 169:28]
      other_state <= 2'h0; // @[IoControl.scala 169:28]
    end else if (_T) begin // @[Conditional.scala 40:58]
      if (dcache_write_other) begin // @[IoControl.scala 183:31]
        other_state <= 2'h3; // @[IoControl.scala 185:20]
      end else if (dcache_read_other) begin // @[IoControl.scala 178:30]
        other_state <= 2'h2; // @[IoControl.scala 181:20]
      end else begin
        other_state <= _GEN_9;
      end
    end else if (_T_1) begin // @[Conditional.scala 39:67]
      other_state <= 2'h0; // @[IoControl.scala 190:18]
    end else if (_T_2) begin // @[Conditional.scala 39:67]
      other_state <= 2'h0; // @[IoControl.scala 194:18]
    end else begin
      other_state <= _GEN_15;
    end
    if (reset) begin // @[IoControl.scala 498:24]
      uart_buffer_0_data <= 8'h0; // @[IoControl.scala 503:13]
    end else if (uart_enq) begin // @[IoControl.scala 403:17]
      if (3'h0 == tail_idx) begin // @[IoControl.scala 404:31]
        uart_buffer_0_data <= io_rxd_uart_data; // @[IoControl.scala 404:31]
      end
    end
    if (reset) begin // @[IoControl.scala 498:24]
      uart_buffer_0_rob_idx <= 3'h0; // @[IoControl.scala 502:16]
    end else if (_GEN_677 == io_rob_commit_1_bits_des_rob & io_rob_commit_1_valid & _GEN_685) begin // @[IoControl.scala 420:138]
      if (3'h0 == flush_head_idx_1) begin // @[IoControl.scala 421:44]
        uart_buffer_0_rob_idx <= 3'h0; // @[IoControl.scala 421:44]
      end else begin
        uart_buffer_0_rob_idx <= _GEN_702;
      end
    end else begin
      uart_buffer_0_rob_idx <= _GEN_702;
    end
    if (reset) begin // @[IoControl.scala 498:24]
      uart_buffer_1_data <= 8'h0; // @[IoControl.scala 503:13]
    end else if (uart_enq) begin // @[IoControl.scala 403:17]
      if (3'h1 == tail_idx) begin // @[IoControl.scala 404:31]
        uart_buffer_1_data <= io_rxd_uart_data; // @[IoControl.scala 404:31]
      end
    end
    if (reset) begin // @[IoControl.scala 498:24]
      uart_buffer_1_rob_idx <= 3'h0; // @[IoControl.scala 502:16]
    end else if (_GEN_677 == io_rob_commit_1_bits_des_rob & io_rob_commit_1_valid & _GEN_685) begin // @[IoControl.scala 420:138]
      if (3'h1 == flush_head_idx_1) begin // @[IoControl.scala 421:44]
        uart_buffer_1_rob_idx <= 3'h0; // @[IoControl.scala 421:44]
      end else begin
        uart_buffer_1_rob_idx <= _GEN_703;
      end
    end else begin
      uart_buffer_1_rob_idx <= _GEN_703;
    end
    if (reset) begin // @[IoControl.scala 498:24]
      uart_buffer_2_data <= 8'h0; // @[IoControl.scala 503:13]
    end else if (uart_enq) begin // @[IoControl.scala 403:17]
      if (3'h2 == tail_idx) begin // @[IoControl.scala 404:31]
        uart_buffer_2_data <= io_rxd_uart_data; // @[IoControl.scala 404:31]
      end
    end
    if (reset) begin // @[IoControl.scala 498:24]
      uart_buffer_2_rob_idx <= 3'h0; // @[IoControl.scala 502:16]
    end else if (_GEN_677 == io_rob_commit_1_bits_des_rob & io_rob_commit_1_valid & _GEN_685) begin // @[IoControl.scala 420:138]
      if (3'h2 == flush_head_idx_1) begin // @[IoControl.scala 421:44]
        uart_buffer_2_rob_idx <= 3'h0; // @[IoControl.scala 421:44]
      end else begin
        uart_buffer_2_rob_idx <= _GEN_704;
      end
    end else begin
      uart_buffer_2_rob_idx <= _GEN_704;
    end
    if (reset) begin // @[IoControl.scala 498:24]
      uart_buffer_3_data <= 8'h0; // @[IoControl.scala 503:13]
    end else if (uart_enq) begin // @[IoControl.scala 403:17]
      if (3'h3 == tail_idx) begin // @[IoControl.scala 404:31]
        uart_buffer_3_data <= io_rxd_uart_data; // @[IoControl.scala 404:31]
      end
    end
    if (reset) begin // @[IoControl.scala 498:24]
      uart_buffer_3_rob_idx <= 3'h0; // @[IoControl.scala 502:16]
    end else if (_GEN_677 == io_rob_commit_1_bits_des_rob & io_rob_commit_1_valid & _GEN_685) begin // @[IoControl.scala 420:138]
      if (3'h3 == flush_head_idx_1) begin // @[IoControl.scala 421:44]
        uart_buffer_3_rob_idx <= 3'h0; // @[IoControl.scala 421:44]
      end else begin
        uart_buffer_3_rob_idx <= _GEN_705;
      end
    end else begin
      uart_buffer_3_rob_idx <= _GEN_705;
    end
    if (reset) begin // @[IoControl.scala 498:24]
      uart_buffer_4_data <= 8'h0; // @[IoControl.scala 503:13]
    end else if (uart_enq) begin // @[IoControl.scala 403:17]
      if (3'h4 == tail_idx) begin // @[IoControl.scala 404:31]
        uart_buffer_4_data <= io_rxd_uart_data; // @[IoControl.scala 404:31]
      end
    end
    if (reset) begin // @[IoControl.scala 498:24]
      uart_buffer_4_rob_idx <= 3'h0; // @[IoControl.scala 502:16]
    end else if (_GEN_677 == io_rob_commit_1_bits_des_rob & io_rob_commit_1_valid & _GEN_685) begin // @[IoControl.scala 420:138]
      if (3'h4 == flush_head_idx_1) begin // @[IoControl.scala 421:44]
        uart_buffer_4_rob_idx <= 3'h0; // @[IoControl.scala 421:44]
      end else begin
        uart_buffer_4_rob_idx <= _GEN_706;
      end
    end else begin
      uart_buffer_4_rob_idx <= _GEN_706;
    end
    if (reset) begin // @[IoControl.scala 498:24]
      uart_buffer_5_data <= 8'h0; // @[IoControl.scala 503:13]
    end else if (uart_enq) begin // @[IoControl.scala 403:17]
      if (3'h5 == tail_idx) begin // @[IoControl.scala 404:31]
        uart_buffer_5_data <= io_rxd_uart_data; // @[IoControl.scala 404:31]
      end
    end
    if (reset) begin // @[IoControl.scala 498:24]
      uart_buffer_5_rob_idx <= 3'h0; // @[IoControl.scala 502:16]
    end else if (_GEN_677 == io_rob_commit_1_bits_des_rob & io_rob_commit_1_valid & _GEN_685) begin // @[IoControl.scala 420:138]
      if (3'h5 == flush_head_idx_1) begin // @[IoControl.scala 421:44]
        uart_buffer_5_rob_idx <= 3'h0; // @[IoControl.scala 421:44]
      end else begin
        uart_buffer_5_rob_idx <= _GEN_707;
      end
    end else begin
      uart_buffer_5_rob_idx <= _GEN_707;
    end
    if (reset) begin // @[IoControl.scala 498:24]
      uart_buffer_6_data <= 8'h0; // @[IoControl.scala 503:13]
    end else if (uart_enq) begin // @[IoControl.scala 403:17]
      if (3'h6 == tail_idx) begin // @[IoControl.scala 404:31]
        uart_buffer_6_data <= io_rxd_uart_data; // @[IoControl.scala 404:31]
      end
    end
    if (reset) begin // @[IoControl.scala 498:24]
      uart_buffer_6_rob_idx <= 3'h0; // @[IoControl.scala 502:16]
    end else if (_GEN_677 == io_rob_commit_1_bits_des_rob & io_rob_commit_1_valid & _GEN_685) begin // @[IoControl.scala 420:138]
      if (3'h6 == flush_head_idx_1) begin // @[IoControl.scala 421:44]
        uart_buffer_6_rob_idx <= 3'h0; // @[IoControl.scala 421:44]
      end else begin
        uart_buffer_6_rob_idx <= _GEN_708;
      end
    end else begin
      uart_buffer_6_rob_idx <= _GEN_708;
    end
    if (reset) begin // @[IoControl.scala 498:24]
      uart_buffer_7_data <= 8'h0; // @[IoControl.scala 503:13]
    end else if (uart_enq) begin // @[IoControl.scala 403:17]
      if (3'h7 == tail_idx) begin // @[IoControl.scala 404:31]
        uart_buffer_7_data <= io_rxd_uart_data; // @[IoControl.scala 404:31]
      end
    end
    if (reset) begin // @[IoControl.scala 498:24]
      uart_buffer_7_rob_idx <= 3'h0; // @[IoControl.scala 502:16]
    end else if (_GEN_677 == io_rob_commit_1_bits_des_rob & io_rob_commit_1_valid & _GEN_685) begin // @[IoControl.scala 420:138]
      if (3'h7 == flush_head_idx_1) begin // @[IoControl.scala 421:44]
        uart_buffer_7_rob_idx <= 3'h0; // @[IoControl.scala 421:44]
      end else begin
        uart_buffer_7_rob_idx <= _GEN_709;
      end
    end else begin
      uart_buffer_7_rob_idx <= _GEN_709;
    end
    if (reset) begin // @[IoControl.scala 379:33]
      uart_buffer_wait_0 <= 1'h0; // @[IoControl.scala 379:33]
    end else if (io_need_flush) begin // @[IoControl.scala 441:22]
      uart_buffer_wait_0 <= 1'h0; // @[IoControl.scala 444:26]
    end else if (_GEN_677 == io_rob_commit_1_bits_des_rob & io_rob_commit_1_valid & _GEN_685) begin // @[IoControl.scala 420:138]
      if (3'h0 == flush_head_idx_1) begin // @[IoControl.scala 422:41]
        uart_buffer_wait_0 <= 1'h0; // @[IoControl.scala 422:41]
      end else begin
        uart_buffer_wait_0 <= _GEN_710;
      end
    end else begin
      uart_buffer_wait_0 <= _GEN_710;
    end
    if (reset) begin // @[IoControl.scala 379:33]
      uart_buffer_wait_1 <= 1'h0; // @[IoControl.scala 379:33]
    end else if (io_need_flush) begin // @[IoControl.scala 441:22]
      uart_buffer_wait_1 <= 1'h0; // @[IoControl.scala 444:26]
    end else if (_GEN_677 == io_rob_commit_1_bits_des_rob & io_rob_commit_1_valid & _GEN_685) begin // @[IoControl.scala 420:138]
      if (3'h1 == flush_head_idx_1) begin // @[IoControl.scala 422:41]
        uart_buffer_wait_1 <= 1'h0; // @[IoControl.scala 422:41]
      end else begin
        uart_buffer_wait_1 <= _GEN_711;
      end
    end else begin
      uart_buffer_wait_1 <= _GEN_711;
    end
    if (reset) begin // @[IoControl.scala 379:33]
      uart_buffer_wait_2 <= 1'h0; // @[IoControl.scala 379:33]
    end else if (io_need_flush) begin // @[IoControl.scala 441:22]
      uart_buffer_wait_2 <= 1'h0; // @[IoControl.scala 444:26]
    end else if (_GEN_677 == io_rob_commit_1_bits_des_rob & io_rob_commit_1_valid & _GEN_685) begin // @[IoControl.scala 420:138]
      if (3'h2 == flush_head_idx_1) begin // @[IoControl.scala 422:41]
        uart_buffer_wait_2 <= 1'h0; // @[IoControl.scala 422:41]
      end else begin
        uart_buffer_wait_2 <= _GEN_712;
      end
    end else begin
      uart_buffer_wait_2 <= _GEN_712;
    end
    if (reset) begin // @[IoControl.scala 379:33]
      uart_buffer_wait_3 <= 1'h0; // @[IoControl.scala 379:33]
    end else if (io_need_flush) begin // @[IoControl.scala 441:22]
      uart_buffer_wait_3 <= 1'h0; // @[IoControl.scala 444:26]
    end else if (_GEN_677 == io_rob_commit_1_bits_des_rob & io_rob_commit_1_valid & _GEN_685) begin // @[IoControl.scala 420:138]
      if (3'h3 == flush_head_idx_1) begin // @[IoControl.scala 422:41]
        uart_buffer_wait_3 <= 1'h0; // @[IoControl.scala 422:41]
      end else begin
        uart_buffer_wait_3 <= _GEN_713;
      end
    end else begin
      uart_buffer_wait_3 <= _GEN_713;
    end
    if (reset) begin // @[IoControl.scala 379:33]
      uart_buffer_wait_4 <= 1'h0; // @[IoControl.scala 379:33]
    end else if (io_need_flush) begin // @[IoControl.scala 441:22]
      uart_buffer_wait_4 <= 1'h0; // @[IoControl.scala 444:26]
    end else if (_GEN_677 == io_rob_commit_1_bits_des_rob & io_rob_commit_1_valid & _GEN_685) begin // @[IoControl.scala 420:138]
      if (3'h4 == flush_head_idx_1) begin // @[IoControl.scala 422:41]
        uart_buffer_wait_4 <= 1'h0; // @[IoControl.scala 422:41]
      end else begin
        uart_buffer_wait_4 <= _GEN_714;
      end
    end else begin
      uart_buffer_wait_4 <= _GEN_714;
    end
    if (reset) begin // @[IoControl.scala 379:33]
      uart_buffer_wait_5 <= 1'h0; // @[IoControl.scala 379:33]
    end else if (io_need_flush) begin // @[IoControl.scala 441:22]
      uart_buffer_wait_5 <= 1'h0; // @[IoControl.scala 444:26]
    end else if (_GEN_677 == io_rob_commit_1_bits_des_rob & io_rob_commit_1_valid & _GEN_685) begin // @[IoControl.scala 420:138]
      if (3'h5 == flush_head_idx_1) begin // @[IoControl.scala 422:41]
        uart_buffer_wait_5 <= 1'h0; // @[IoControl.scala 422:41]
      end else begin
        uart_buffer_wait_5 <= _GEN_715;
      end
    end else begin
      uart_buffer_wait_5 <= _GEN_715;
    end
    if (reset) begin // @[IoControl.scala 379:33]
      uart_buffer_wait_6 <= 1'h0; // @[IoControl.scala 379:33]
    end else if (io_need_flush) begin // @[IoControl.scala 441:22]
      uart_buffer_wait_6 <= 1'h0; // @[IoControl.scala 444:26]
    end else if (_GEN_677 == io_rob_commit_1_bits_des_rob & io_rob_commit_1_valid & _GEN_685) begin // @[IoControl.scala 420:138]
      if (3'h6 == flush_head_idx_1) begin // @[IoControl.scala 422:41]
        uart_buffer_wait_6 <= 1'h0; // @[IoControl.scala 422:41]
      end else begin
        uart_buffer_wait_6 <= _GEN_716;
      end
    end else begin
      uart_buffer_wait_6 <= _GEN_716;
    end
    if (reset) begin // @[IoControl.scala 379:33]
      uart_buffer_wait_7 <= 1'h0; // @[IoControl.scala 379:33]
    end else if (io_need_flush) begin // @[IoControl.scala 441:22]
      uart_buffer_wait_7 <= 1'h0; // @[IoControl.scala 444:26]
    end else if (_GEN_677 == io_rob_commit_1_bits_des_rob & io_rob_commit_1_valid & _GEN_685) begin // @[IoControl.scala 420:138]
      if (3'h7 == flush_head_idx_1) begin // @[IoControl.scala 422:41]
        uart_buffer_wait_7 <= 1'h0; // @[IoControl.scala 422:41]
      end else begin
        uart_buffer_wait_7 <= _GEN_717;
      end
    end else begin
      uart_buffer_wait_7 <= _GEN_717;
    end
    if (reset) begin // @[IoControl.scala 380:26]
      uart_head <= 8'h1; // @[IoControl.scala 380:26]
    end else if (io_need_flush) begin // @[IoControl.scala 441:22]
      if (will_drop_1) begin // @[IoControl.scala 427:84]
        uart_head <= _next_flush_head_T_2;
      end else if (will_drop_0) begin // @[IoControl.scala 427:84]
        uart_head <= _flush_head_idx_T_2;
      end else begin
        uart_head <= uart_flush_head;
      end
    end else if (uart_deq) begin // @[IoControl.scala 409:18]
      uart_head <= _uart_head_T; // @[IoControl.scala 412:14]
    end
    if (reset) begin // @[IoControl.scala 382:32]
      uart_flush_head <= 8'h1; // @[IoControl.scala 382:32]
    end else if (will_drop_1) begin // @[IoControl.scala 427:84]
      uart_flush_head <= _next_flush_head_T_2;
    end else if (will_drop_0) begin // @[IoControl.scala 427:84]
      uart_flush_head <= _flush_head_idx_T_2;
    end
    if (reset) begin // @[IoControl.scala 383:26]
      uart_tail <= 8'h1; // @[IoControl.scala 383:26]
    end else if (uart_enq) begin // @[IoControl.scala 403:17]
      uart_tail <= _uart_tail_T; // @[IoControl.scala 406:14]
    end
    if (reset) begin // @[IoControl.scala 385:27]
      maybe_full <= 1'h0; // @[IoControl.scala 385:27]
    end else if (io_need_flush) begin // @[IoControl.scala 441:22]
      maybe_full <= maybe_true_full; // @[IoControl.scala 446:15]
    end else begin
      maybe_full <= _GEN_755;
    end
    if (reset) begin // @[IoControl.scala 386:32]
      maybe_true_full <= 1'h0; // @[IoControl.scala 386:32]
    end else begin
      maybe_true_full <= _GEN_753;
    end
    if (reset) begin // @[IoControl.scala 452:27]
      uart_state <= 2'h0; // @[IoControl.scala 452:27]
    end else if (_T_56) begin // @[Conditional.scala 40:58]
      if (dcache_write_uart & ~io_txd_uart_busy) begin // @[IoControl.scala 470:50]
        uart_state <= 2'h2; // @[IoControl.scala 474:19]
      end else if (dcache_read_uart & _uart_deq_T) begin // @[IoControl.scala 475:48]
        uart_state <= 2'h1; // @[IoControl.scala 480:19]
      end else begin
        uart_state <= _GEN_770;
      end
    end else if (_T_60) begin // @[Conditional.scala 39:67]
      uart_state <= 2'h0; // @[IoControl.scala 489:17]
    end else if (_T_61) begin // @[Conditional.scala 39:67]
      uart_state <= 2'h0; // @[IoControl.scala 493:17]
    end
    if (reset) begin // @[IoControl.scala 453:31]
      txd_uart_start <= 1'h0; // @[IoControl.scala 453:31]
    end else if (_T_56) begin // @[Conditional.scala 40:58]
      txd_uart_start <= _GEN_776;
    end else if (_T_60) begin // @[Conditional.scala 39:67]
      txd_uart_start <= 1'h0; // @[IoControl.scala 488:21]
    end
    if (reset) begin // @[IoControl.scala 454:30]
      txd_uart_data <= 8'h0; // @[IoControl.scala 454:30]
    end else if (_T_56) begin // @[Conditional.scala 40:58]
      if (dcache_write_uart & ~io_txd_uart_busy) begin // @[IoControl.scala 470:50]
        txd_uart_data <= io_dcache_write_req_bits_data[7:0]; // @[IoControl.scala 472:22]
      end
    end
  end
// Register and memory initialization
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  base_ram_ctrl_data_out = _RAND_0[31:0];
  _RAND_1 = {1{`RANDOM}};
  base_ram_ctrl_addr = _RAND_1[19:0];
  _RAND_2 = {1{`RANDOM}};
  base_ram_ctrl_be_n = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  base_ram_ctrl_ce_n = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  base_ram_ctrl_oe_n = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  base_ram_ctrl_we_n = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  ext_ram_ctrl_data_out = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  ext_ram_ctrl_addr = _RAND_7[19:0];
  _RAND_8 = {1{`RANDOM}};
  ext_ram_ctrl_be_n = _RAND_8[3:0];
  _RAND_9 = {1{`RANDOM}};
  ext_ram_ctrl_ce_n = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  ext_ram_ctrl_oe_n = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  ext_ram_ctrl_we_n = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  base_state = _RAND_12[2:0];
  _RAND_13 = {1{`RANDOM}};
  base_clock_counter = _RAND_13[3:0];
  _RAND_14 = {1{`RANDOM}};
  base_wait_counter = _RAND_14[3:0];
  _RAND_15 = {1{`RANDOM}};
  ext_state = _RAND_15[2:0];
  _RAND_16 = {1{`RANDOM}};
  ext_clock_counter = _RAND_16[3:0];
  _RAND_17 = {1{`RANDOM}};
  ext_wait_counter = _RAND_17[3:0];
  _RAND_18 = {1{`RANDOM}};
  icache_buffer_0 = _RAND_18[31:0];
  _RAND_19 = {1{`RANDOM}};
  icache_buffer_1 = _RAND_19[31:0];
  _RAND_20 = {1{`RANDOM}};
  icache_buffer_2 = _RAND_20[31:0];
  _RAND_21 = {1{`RANDOM}};
  icache_buffer_3 = _RAND_21[31:0];
  _RAND_22 = {1{`RANDOM}};
  icache_buffer_4 = _RAND_22[31:0];
  _RAND_23 = {1{`RANDOM}};
  icache_buffer_5 = _RAND_23[31:0];
  _RAND_24 = {1{`RANDOM}};
  icache_buffer_6 = _RAND_24[31:0];
  _RAND_25 = {1{`RANDOM}};
  icache_buffer_7 = _RAND_25[31:0];
  _RAND_26 = {1{`RANDOM}};
  icache_data_valid = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  dcache_buffer = _RAND_27[31:0];
  _RAND_28 = {1{`RANDOM}};
  dcache_data_valid = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  other_state = _RAND_29[1:0];
  _RAND_30 = {1{`RANDOM}};
  uart_buffer_0_data = _RAND_30[7:0];
  _RAND_31 = {1{`RANDOM}};
  uart_buffer_0_rob_idx = _RAND_31[2:0];
  _RAND_32 = {1{`RANDOM}};
  uart_buffer_1_data = _RAND_32[7:0];
  _RAND_33 = {1{`RANDOM}};
  uart_buffer_1_rob_idx = _RAND_33[2:0];
  _RAND_34 = {1{`RANDOM}};
  uart_buffer_2_data = _RAND_34[7:0];
  _RAND_35 = {1{`RANDOM}};
  uart_buffer_2_rob_idx = _RAND_35[2:0];
  _RAND_36 = {1{`RANDOM}};
  uart_buffer_3_data = _RAND_36[7:0];
  _RAND_37 = {1{`RANDOM}};
  uart_buffer_3_rob_idx = _RAND_37[2:0];
  _RAND_38 = {1{`RANDOM}};
  uart_buffer_4_data = _RAND_38[7:0];
  _RAND_39 = {1{`RANDOM}};
  uart_buffer_4_rob_idx = _RAND_39[2:0];
  _RAND_40 = {1{`RANDOM}};
  uart_buffer_5_data = _RAND_40[7:0];
  _RAND_41 = {1{`RANDOM}};
  uart_buffer_5_rob_idx = _RAND_41[2:0];
  _RAND_42 = {1{`RANDOM}};
  uart_buffer_6_data = _RAND_42[7:0];
  _RAND_43 = {1{`RANDOM}};
  uart_buffer_6_rob_idx = _RAND_43[2:0];
  _RAND_44 = {1{`RANDOM}};
  uart_buffer_7_data = _RAND_44[7:0];
  _RAND_45 = {1{`RANDOM}};
  uart_buffer_7_rob_idx = _RAND_45[2:0];
  _RAND_46 = {1{`RANDOM}};
  uart_buffer_wait_0 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  uart_buffer_wait_1 = _RAND_47[0:0];
  _RAND_48 = {1{`RANDOM}};
  uart_buffer_wait_2 = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  uart_buffer_wait_3 = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  uart_buffer_wait_4 = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  uart_buffer_wait_5 = _RAND_51[0:0];
  _RAND_52 = {1{`RANDOM}};
  uart_buffer_wait_6 = _RAND_52[0:0];
  _RAND_53 = {1{`RANDOM}};
  uart_buffer_wait_7 = _RAND_53[0:0];
  _RAND_54 = {1{`RANDOM}};
  uart_head = _RAND_54[7:0];
  _RAND_55 = {1{`RANDOM}};
  uart_flush_head = _RAND_55[7:0];
  _RAND_56 = {1{`RANDOM}};
  uart_tail = _RAND_56[7:0];
  _RAND_57 = {1{`RANDOM}};
  maybe_full = _RAND_57[0:0];
  _RAND_58 = {1{`RANDOM}};
  maybe_true_full = _RAND_58[0:0];
  _RAND_59 = {1{`RANDOM}};
  uart_state = _RAND_59[1:0];
  _RAND_60 = {1{`RANDOM}};
  txd_uart_start = _RAND_60[0:0];
  _RAND_61 = {1{`RANDOM}};
  txd_uart_data = _RAND_61[7:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
endmodule
module Top(
  input         clock,
  input         reset,
  input  [31:0] io_base_ram_ctrl_data_in,
  output [31:0] io_base_ram_ctrl_ctrl_data_out,
  output [19:0] io_base_ram_ctrl_ctrl_addr,
  output [3:0]  io_base_ram_ctrl_ctrl_be_n,
  output        io_base_ram_ctrl_ctrl_ce_n,
  output        io_base_ram_ctrl_ctrl_oe_n,
  output        io_base_ram_ctrl_ctrl_we_n,
  input  [31:0] io_ext_ram_ctrl_data_in,
  output [31:0] io_ext_ram_ctrl_ctrl_data_out,
  output [19:0] io_ext_ram_ctrl_ctrl_addr,
  output [3:0]  io_ext_ram_ctrl_ctrl_be_n,
  output        io_ext_ram_ctrl_ctrl_ce_n,
  output        io_ext_ram_ctrl_ctrl_oe_n,
  output        io_ext_ram_ctrl_ctrl_we_n,
  input         io_rxd_uart_ready,
  output        io_rxd_uart_clear,
  input  [7:0]  io_rxd_uart_data,
  output        io_txd_uart_start,
  output [7:0]  io_txd_uart_data,
  input         io_txd_uart_busy,
  output [2:0]  io_io_control_debug_base_state,
  output        io_io_control_debug_icache_read_base,
  output        io_io_control_debug_icache_read_ext,
  output        io_io_control_debug_dcache_read_base,
  output        io_io_control_debug_dcache_read_ext,
  output        io_io_control_debug_dcache_write_base,
  output        io_io_control_debug_dcache_write_ext,
  output [19:0] io_io_control_debug_icache_read_addr,
  output [19:0] io_io_control_debug_dcache_read_addr,
  output [19:0] io_io_control_debug_dcache_write_addr,
  output        io_icache_debug_state,
  output        io_icache_debug_hit_cache,
  output        io_icache_debug_cache_we,
  output [19:0] io_icache_debug_cache_read_tag,
  output        io_icache_debug_icache_req_valid,
  output [31:0] io_icache_debug_icache_req_bits_addr,
  output [7:0]  io_bpu_debug_branch_mask,
  output [7:0]  io_bpu_debug_fetched_mask,
  output [7:0]  io_bpu_debug_predict_branch,
  output [31:0] io_bpu_debug_predict_addr,
  output        io_bpu_debug_is_taken,
  output        io_bpu_debug_take_delay,
  output [31:0] io_bpu_debug_inst_packet_0,
  output [31:0] io_bpu_debug_inst_packet_1,
  output [31:0] io_bpu_debug_inst_packet_2,
  output [31:0] io_bpu_debug_inst_packet_3,
  output [31:0] io_bpu_debug_inst_packet_4,
  output [31:0] io_bpu_debug_inst_packet_5,
  output [31:0] io_bpu_debug_inst_packet_6,
  output [31:0] io_bpu_debug_inst_packet_7
);
  wire  core_clock; // @[Top.scala 17:20]
  wire  core_reset; // @[Top.scala 17:20]
  wire  core_io_icache_io_read_req_ready; // @[Top.scala 17:20]
  wire  core_io_icache_io_read_req_valid; // @[Top.scala 17:20]
  wire [31:0] core_io_icache_io_read_req_bits_addr; // @[Top.scala 17:20]
  wire [255:0] core_io_icache_io_read_resp_bits_data; // @[Top.scala 17:20]
  wire  core_io_dcache_io_read_req_ready; // @[Top.scala 17:20]
  wire  core_io_dcache_io_read_req_valid; // @[Top.scala 17:20]
  wire [31:0] core_io_dcache_io_read_req_bits_addr; // @[Top.scala 17:20]
  wire [3:0] core_io_dcache_io_read_req_bits_rob_idx; // @[Top.scala 17:20]
  wire [31:0] core_io_dcache_io_read_resp_bits_data; // @[Top.scala 17:20]
  wire  core_io_dcache_io_write_req_ready; // @[Top.scala 17:20]
  wire  core_io_dcache_io_write_req_valid; // @[Top.scala 17:20]
  wire [31:0] core_io_dcache_io_write_req_bits_addr; // @[Top.scala 17:20]
  wire [31:0] core_io_dcache_io_write_req_bits_data; // @[Top.scala 17:20]
  wire [3:0] core_io_dcache_io_write_req_bits_byte_mask; // @[Top.scala 17:20]
  wire  core_io_need_flush; // @[Top.scala 17:20]
  wire  core_io_rob_commit_0_valid; // @[Top.scala 17:20]
  wire [2:0] core_io_rob_commit_0_bits_des_rob; // @[Top.scala 17:20]
  wire  core_io_rob_commit_1_valid; // @[Top.scala 17:20]
  wire [2:0] core_io_rob_commit_1_bits_des_rob; // @[Top.scala 17:20]
  wire  core_io_icache_debug_state; // @[Top.scala 17:20]
  wire  core_io_icache_debug_hit_cache; // @[Top.scala 17:20]
  wire  core_io_icache_debug_cache_we; // @[Top.scala 17:20]
  wire [19:0] core_io_icache_debug_cache_read_tag; // @[Top.scala 17:20]
  wire  core_io_icache_debug_icache_req_valid; // @[Top.scala 17:20]
  wire [31:0] core_io_icache_debug_icache_req_bits_addr; // @[Top.scala 17:20]
  wire [7:0] core_io_bpu_debug_branch_mask; // @[Top.scala 17:20]
  wire [7:0] core_io_bpu_debug_fetched_mask; // @[Top.scala 17:20]
  wire [7:0] core_io_bpu_debug_predict_branch; // @[Top.scala 17:20]
  wire [31:0] core_io_bpu_debug_predict_addr; // @[Top.scala 17:20]
  wire  core_io_bpu_debug_is_taken; // @[Top.scala 17:20]
  wire  core_io_bpu_debug_take_delay; // @[Top.scala 17:20]
  wire [31:0] core_io_bpu_debug_inst_packet_0; // @[Top.scala 17:20]
  wire [31:0] core_io_bpu_debug_inst_packet_1; // @[Top.scala 17:20]
  wire [31:0] core_io_bpu_debug_inst_packet_2; // @[Top.scala 17:20]
  wire [31:0] core_io_bpu_debug_inst_packet_3; // @[Top.scala 17:20]
  wire [31:0] core_io_bpu_debug_inst_packet_4; // @[Top.scala 17:20]
  wire [31:0] core_io_bpu_debug_inst_packet_5; // @[Top.scala 17:20]
  wire [31:0] core_io_bpu_debug_inst_packet_6; // @[Top.scala 17:20]
  wire [31:0] core_io_bpu_debug_inst_packet_7; // @[Top.scala 17:20]
  wire  io_control_clock; // @[Top.scala 18:26]
  wire  io_control_reset; // @[Top.scala 18:26]
  wire  io_control_io_icache_read_req_ready; // @[Top.scala 18:26]
  wire  io_control_io_icache_read_req_valid; // @[Top.scala 18:26]
  wire [31:0] io_control_io_icache_read_req_bits_addr; // @[Top.scala 18:26]
  wire [255:0] io_control_io_icache_read_resp_bits_data; // @[Top.scala 18:26]
  wire  io_control_io_dcache_read_req_ready; // @[Top.scala 18:26]
  wire  io_control_io_dcache_read_req_valid; // @[Top.scala 18:26]
  wire [31:0] io_control_io_dcache_read_req_bits_addr; // @[Top.scala 18:26]
  wire [3:0] io_control_io_dcache_read_req_bits_rob_idx; // @[Top.scala 18:26]
  wire [31:0] io_control_io_dcache_read_resp_bits_data; // @[Top.scala 18:26]
  wire  io_control_io_dcache_write_req_ready; // @[Top.scala 18:26]
  wire  io_control_io_dcache_write_req_valid; // @[Top.scala 18:26]
  wire [31:0] io_control_io_dcache_write_req_bits_addr; // @[Top.scala 18:26]
  wire [31:0] io_control_io_dcache_write_req_bits_data; // @[Top.scala 18:26]
  wire [3:0] io_control_io_dcache_write_req_bits_byte_mask; // @[Top.scala 18:26]
  wire [31:0] io_control_io_base_ram_ctrl_data_in; // @[Top.scala 18:26]
  wire [31:0] io_control_io_base_ram_ctrl_ctrl_data_out; // @[Top.scala 18:26]
  wire [19:0] io_control_io_base_ram_ctrl_ctrl_addr; // @[Top.scala 18:26]
  wire [3:0] io_control_io_base_ram_ctrl_ctrl_be_n; // @[Top.scala 18:26]
  wire  io_control_io_base_ram_ctrl_ctrl_ce_n; // @[Top.scala 18:26]
  wire  io_control_io_base_ram_ctrl_ctrl_oe_n; // @[Top.scala 18:26]
  wire  io_control_io_base_ram_ctrl_ctrl_we_n; // @[Top.scala 18:26]
  wire [31:0] io_control_io_ext_ram_ctrl_data_in; // @[Top.scala 18:26]
  wire [31:0] io_control_io_ext_ram_ctrl_ctrl_data_out; // @[Top.scala 18:26]
  wire [19:0] io_control_io_ext_ram_ctrl_ctrl_addr; // @[Top.scala 18:26]
  wire [3:0] io_control_io_ext_ram_ctrl_ctrl_be_n; // @[Top.scala 18:26]
  wire  io_control_io_ext_ram_ctrl_ctrl_ce_n; // @[Top.scala 18:26]
  wire  io_control_io_ext_ram_ctrl_ctrl_oe_n; // @[Top.scala 18:26]
  wire  io_control_io_ext_ram_ctrl_ctrl_we_n; // @[Top.scala 18:26]
  wire  io_control_io_rxd_uart_ready; // @[Top.scala 18:26]
  wire  io_control_io_rxd_uart_clear; // @[Top.scala 18:26]
  wire [7:0] io_control_io_rxd_uart_data; // @[Top.scala 18:26]
  wire  io_control_io_txd_uart_start; // @[Top.scala 18:26]
  wire [7:0] io_control_io_txd_uart_data; // @[Top.scala 18:26]
  wire  io_control_io_txd_uart_busy; // @[Top.scala 18:26]
  wire  io_control_io_rob_commit_0_valid; // @[Top.scala 18:26]
  wire [2:0] io_control_io_rob_commit_0_bits_des_rob; // @[Top.scala 18:26]
  wire  io_control_io_rob_commit_1_valid; // @[Top.scala 18:26]
  wire [2:0] io_control_io_rob_commit_1_bits_des_rob; // @[Top.scala 18:26]
  wire  io_control_io_need_flush; // @[Top.scala 18:26]
  wire [2:0] io_control_io_debug_base_state; // @[Top.scala 18:26]
  wire  io_control_io_debug_icache_read_base; // @[Top.scala 18:26]
  wire  io_control_io_debug_icache_read_ext; // @[Top.scala 18:26]
  wire  io_control_io_debug_dcache_read_base; // @[Top.scala 18:26]
  wire  io_control_io_debug_dcache_read_ext; // @[Top.scala 18:26]
  wire  io_control_io_debug_dcache_write_base; // @[Top.scala 18:26]
  wire  io_control_io_debug_dcache_write_ext; // @[Top.scala 18:26]
  wire [19:0] io_control_io_debug_icache_read_addr; // @[Top.scala 18:26]
  wire [19:0] io_control_io_debug_dcache_read_addr; // @[Top.scala 18:26]
  wire [19:0] io_control_io_debug_dcache_write_addr; // @[Top.scala 18:26]
  Core core ( // @[Top.scala 17:20]
    .clock(core_clock),
    .reset(core_reset),
    .io_icache_io_read_req_ready(core_io_icache_io_read_req_ready),
    .io_icache_io_read_req_valid(core_io_icache_io_read_req_valid),
    .io_icache_io_read_req_bits_addr(core_io_icache_io_read_req_bits_addr),
    .io_icache_io_read_resp_bits_data(core_io_icache_io_read_resp_bits_data),
    .io_dcache_io_read_req_ready(core_io_dcache_io_read_req_ready),
    .io_dcache_io_read_req_valid(core_io_dcache_io_read_req_valid),
    .io_dcache_io_read_req_bits_addr(core_io_dcache_io_read_req_bits_addr),
    .io_dcache_io_read_req_bits_rob_idx(core_io_dcache_io_read_req_bits_rob_idx),
    .io_dcache_io_read_resp_bits_data(core_io_dcache_io_read_resp_bits_data),
    .io_dcache_io_write_req_ready(core_io_dcache_io_write_req_ready),
    .io_dcache_io_write_req_valid(core_io_dcache_io_write_req_valid),
    .io_dcache_io_write_req_bits_addr(core_io_dcache_io_write_req_bits_addr),
    .io_dcache_io_write_req_bits_data(core_io_dcache_io_write_req_bits_data),
    .io_dcache_io_write_req_bits_byte_mask(core_io_dcache_io_write_req_bits_byte_mask),
    .io_need_flush(core_io_need_flush),
    .io_rob_commit_0_valid(core_io_rob_commit_0_valid),
    .io_rob_commit_0_bits_des_rob(core_io_rob_commit_0_bits_des_rob),
    .io_rob_commit_1_valid(core_io_rob_commit_1_valid),
    .io_rob_commit_1_bits_des_rob(core_io_rob_commit_1_bits_des_rob),
    .io_icache_debug_state(core_io_icache_debug_state),
    .io_icache_debug_hit_cache(core_io_icache_debug_hit_cache),
    .io_icache_debug_cache_we(core_io_icache_debug_cache_we),
    .io_icache_debug_cache_read_tag(core_io_icache_debug_cache_read_tag),
    .io_icache_debug_icache_req_valid(core_io_icache_debug_icache_req_valid),
    .io_icache_debug_icache_req_bits_addr(core_io_icache_debug_icache_req_bits_addr),
    .io_bpu_debug_branch_mask(core_io_bpu_debug_branch_mask),
    .io_bpu_debug_fetched_mask(core_io_bpu_debug_fetched_mask),
    .io_bpu_debug_predict_branch(core_io_bpu_debug_predict_branch),
    .io_bpu_debug_predict_addr(core_io_bpu_debug_predict_addr),
    .io_bpu_debug_is_taken(core_io_bpu_debug_is_taken),
    .io_bpu_debug_take_delay(core_io_bpu_debug_take_delay),
    .io_bpu_debug_inst_packet_0(core_io_bpu_debug_inst_packet_0),
    .io_bpu_debug_inst_packet_1(core_io_bpu_debug_inst_packet_1),
    .io_bpu_debug_inst_packet_2(core_io_bpu_debug_inst_packet_2),
    .io_bpu_debug_inst_packet_3(core_io_bpu_debug_inst_packet_3),
    .io_bpu_debug_inst_packet_4(core_io_bpu_debug_inst_packet_4),
    .io_bpu_debug_inst_packet_5(core_io_bpu_debug_inst_packet_5),
    .io_bpu_debug_inst_packet_6(core_io_bpu_debug_inst_packet_6),
    .io_bpu_debug_inst_packet_7(core_io_bpu_debug_inst_packet_7)
  );
  IoControl io_control ( // @[Top.scala 18:26]
    .clock(io_control_clock),
    .reset(io_control_reset),
    .io_icache_read_req_ready(io_control_io_icache_read_req_ready),
    .io_icache_read_req_valid(io_control_io_icache_read_req_valid),
    .io_icache_read_req_bits_addr(io_control_io_icache_read_req_bits_addr),
    .io_icache_read_resp_bits_data(io_control_io_icache_read_resp_bits_data),
    .io_dcache_read_req_ready(io_control_io_dcache_read_req_ready),
    .io_dcache_read_req_valid(io_control_io_dcache_read_req_valid),
    .io_dcache_read_req_bits_addr(io_control_io_dcache_read_req_bits_addr),
    .io_dcache_read_req_bits_rob_idx(io_control_io_dcache_read_req_bits_rob_idx),
    .io_dcache_read_resp_bits_data(io_control_io_dcache_read_resp_bits_data),
    .io_dcache_write_req_ready(io_control_io_dcache_write_req_ready),
    .io_dcache_write_req_valid(io_control_io_dcache_write_req_valid),
    .io_dcache_write_req_bits_addr(io_control_io_dcache_write_req_bits_addr),
    .io_dcache_write_req_bits_data(io_control_io_dcache_write_req_bits_data),
    .io_dcache_write_req_bits_byte_mask(io_control_io_dcache_write_req_bits_byte_mask),
    .io_base_ram_ctrl_data_in(io_control_io_base_ram_ctrl_data_in),
    .io_base_ram_ctrl_ctrl_data_out(io_control_io_base_ram_ctrl_ctrl_data_out),
    .io_base_ram_ctrl_ctrl_addr(io_control_io_base_ram_ctrl_ctrl_addr),
    .io_base_ram_ctrl_ctrl_be_n(io_control_io_base_ram_ctrl_ctrl_be_n),
    .io_base_ram_ctrl_ctrl_ce_n(io_control_io_base_ram_ctrl_ctrl_ce_n),
    .io_base_ram_ctrl_ctrl_oe_n(io_control_io_base_ram_ctrl_ctrl_oe_n),
    .io_base_ram_ctrl_ctrl_we_n(io_control_io_base_ram_ctrl_ctrl_we_n),
    .io_ext_ram_ctrl_data_in(io_control_io_ext_ram_ctrl_data_in),
    .io_ext_ram_ctrl_ctrl_data_out(io_control_io_ext_ram_ctrl_ctrl_data_out),
    .io_ext_ram_ctrl_ctrl_addr(io_control_io_ext_ram_ctrl_ctrl_addr),
    .io_ext_ram_ctrl_ctrl_be_n(io_control_io_ext_ram_ctrl_ctrl_be_n),
    .io_ext_ram_ctrl_ctrl_ce_n(io_control_io_ext_ram_ctrl_ctrl_ce_n),
    .io_ext_ram_ctrl_ctrl_oe_n(io_control_io_ext_ram_ctrl_ctrl_oe_n),
    .io_ext_ram_ctrl_ctrl_we_n(io_control_io_ext_ram_ctrl_ctrl_we_n),
    .io_rxd_uart_ready(io_control_io_rxd_uart_ready),
    .io_rxd_uart_clear(io_control_io_rxd_uart_clear),
    .io_rxd_uart_data(io_control_io_rxd_uart_data),
    .io_txd_uart_start(io_control_io_txd_uart_start),
    .io_txd_uart_data(io_control_io_txd_uart_data),
    .io_txd_uart_busy(io_control_io_txd_uart_busy),
    .io_rob_commit_0_valid(io_control_io_rob_commit_0_valid),
    .io_rob_commit_0_bits_des_rob(io_control_io_rob_commit_0_bits_des_rob),
    .io_rob_commit_1_valid(io_control_io_rob_commit_1_valid),
    .io_rob_commit_1_bits_des_rob(io_control_io_rob_commit_1_bits_des_rob),
    .io_need_flush(io_control_io_need_flush),
    .io_debug_base_state(io_control_io_debug_base_state),
    .io_debug_icache_read_base(io_control_io_debug_icache_read_base),
    .io_debug_icache_read_ext(io_control_io_debug_icache_read_ext),
    .io_debug_dcache_read_base(io_control_io_debug_dcache_read_base),
    .io_debug_dcache_read_ext(io_control_io_debug_dcache_read_ext),
    .io_debug_dcache_write_base(io_control_io_debug_dcache_write_base),
    .io_debug_dcache_write_ext(io_control_io_debug_dcache_write_ext),
    .io_debug_icache_read_addr(io_control_io_debug_icache_read_addr),
    .io_debug_dcache_read_addr(io_control_io_debug_dcache_read_addr),
    .io_debug_dcache_write_addr(io_control_io_debug_dcache_write_addr)
  );
  assign io_base_ram_ctrl_ctrl_data_out = io_control_io_base_ram_ctrl_ctrl_data_out; // @[Top.scala 28:19]
  assign io_base_ram_ctrl_ctrl_addr = io_control_io_base_ram_ctrl_ctrl_addr; // @[Top.scala 28:19]
  assign io_base_ram_ctrl_ctrl_be_n = io_control_io_base_ram_ctrl_ctrl_be_n; // @[Top.scala 28:19]
  assign io_base_ram_ctrl_ctrl_ce_n = io_control_io_base_ram_ctrl_ctrl_ce_n; // @[Top.scala 28:19]
  assign io_base_ram_ctrl_ctrl_oe_n = io_control_io_base_ram_ctrl_ctrl_oe_n; // @[Top.scala 28:19]
  assign io_base_ram_ctrl_ctrl_we_n = io_control_io_base_ram_ctrl_ctrl_we_n; // @[Top.scala 28:19]
  assign io_ext_ram_ctrl_ctrl_data_out = io_control_io_ext_ram_ctrl_ctrl_data_out; // @[Top.scala 27:18]
  assign io_ext_ram_ctrl_ctrl_addr = io_control_io_ext_ram_ctrl_ctrl_addr; // @[Top.scala 27:18]
  assign io_ext_ram_ctrl_ctrl_be_n = io_control_io_ext_ram_ctrl_ctrl_be_n; // @[Top.scala 27:18]
  assign io_ext_ram_ctrl_ctrl_ce_n = io_control_io_ext_ram_ctrl_ctrl_ce_n; // @[Top.scala 27:18]
  assign io_ext_ram_ctrl_ctrl_oe_n = io_control_io_ext_ram_ctrl_ctrl_oe_n; // @[Top.scala 27:18]
  assign io_ext_ram_ctrl_ctrl_we_n = io_control_io_ext_ram_ctrl_ctrl_we_n; // @[Top.scala 27:18]
  assign io_rxd_uart_clear = io_control_io_rxd_uart_clear; // @[Top.scala 29:9]
  assign io_txd_uart_start = io_control_io_txd_uart_start; // @[Top.scala 30:9]
  assign io_txd_uart_data = io_control_io_txd_uart_data; // @[Top.scala 30:9]
  assign io_io_control_debug_base_state = io_control_io_debug_base_state; // @[Top.scala 32:22]
  assign io_io_control_debug_icache_read_base = io_control_io_debug_icache_read_base; // @[Top.scala 32:22]
  assign io_io_control_debug_icache_read_ext = io_control_io_debug_icache_read_ext; // @[Top.scala 32:22]
  assign io_io_control_debug_dcache_read_base = io_control_io_debug_dcache_read_base; // @[Top.scala 32:22]
  assign io_io_control_debug_dcache_read_ext = io_control_io_debug_dcache_read_ext; // @[Top.scala 32:22]
  assign io_io_control_debug_dcache_write_base = io_control_io_debug_dcache_write_base; // @[Top.scala 32:22]
  assign io_io_control_debug_dcache_write_ext = io_control_io_debug_dcache_write_ext; // @[Top.scala 32:22]
  assign io_io_control_debug_icache_read_addr = io_control_io_debug_icache_read_addr; // @[Top.scala 32:22]
  assign io_io_control_debug_dcache_read_addr = io_control_io_debug_dcache_read_addr; // @[Top.scala 32:22]
  assign io_io_control_debug_dcache_write_addr = io_control_io_debug_dcache_write_addr; // @[Top.scala 32:22]
  assign io_icache_debug_state = core_io_icache_debug_state; // @[Top.scala 33:18]
  assign io_icache_debug_hit_cache = core_io_icache_debug_hit_cache; // @[Top.scala 33:18]
  assign io_icache_debug_cache_we = core_io_icache_debug_cache_we; // @[Top.scala 33:18]
  assign io_icache_debug_cache_read_tag = core_io_icache_debug_cache_read_tag; // @[Top.scala 33:18]
  assign io_icache_debug_icache_req_valid = core_io_icache_debug_icache_req_valid; // @[Top.scala 33:18]
  assign io_icache_debug_icache_req_bits_addr = core_io_icache_debug_icache_req_bits_addr; // @[Top.scala 33:18]
  assign io_bpu_debug_branch_mask = core_io_bpu_debug_branch_mask; // @[Top.scala 34:15]
  assign io_bpu_debug_fetched_mask = core_io_bpu_debug_fetched_mask; // @[Top.scala 34:15]
  assign io_bpu_debug_predict_branch = core_io_bpu_debug_predict_branch; // @[Top.scala 34:15]
  assign io_bpu_debug_predict_addr = core_io_bpu_debug_predict_addr; // @[Top.scala 34:15]
  assign io_bpu_debug_is_taken = core_io_bpu_debug_is_taken; // @[Top.scala 34:15]
  assign io_bpu_debug_take_delay = core_io_bpu_debug_take_delay; // @[Top.scala 34:15]
  assign io_bpu_debug_inst_packet_0 = core_io_bpu_debug_inst_packet_0; // @[Top.scala 34:15]
  assign io_bpu_debug_inst_packet_1 = core_io_bpu_debug_inst_packet_1; // @[Top.scala 34:15]
  assign io_bpu_debug_inst_packet_2 = core_io_bpu_debug_inst_packet_2; // @[Top.scala 34:15]
  assign io_bpu_debug_inst_packet_3 = core_io_bpu_debug_inst_packet_3; // @[Top.scala 34:15]
  assign io_bpu_debug_inst_packet_4 = core_io_bpu_debug_inst_packet_4; // @[Top.scala 34:15]
  assign io_bpu_debug_inst_packet_5 = core_io_bpu_debug_inst_packet_5; // @[Top.scala 34:15]
  assign io_bpu_debug_inst_packet_6 = core_io_bpu_debug_inst_packet_6; // @[Top.scala 34:15]
  assign io_bpu_debug_inst_packet_7 = core_io_bpu_debug_inst_packet_7; // @[Top.scala 34:15]
  assign core_clock = clock;
  assign core_reset = reset;
  assign core_io_icache_io_read_req_ready = io_control_io_icache_read_req_ready; // @[Top.scala 19:30]
  assign core_io_icache_io_read_resp_bits_data = io_control_io_icache_read_resp_bits_data; // @[Top.scala 20:30]
  assign core_io_dcache_io_read_req_ready = io_control_io_dcache_read_req_ready; // @[Top.scala 21:30]
  assign core_io_dcache_io_read_resp_bits_data = io_control_io_dcache_read_resp_bits_data; // @[Top.scala 22:30]
  assign core_io_dcache_io_write_req_ready = io_control_io_dcache_write_req_ready; // @[Top.scala 23:30]
  assign io_control_clock = clock;
  assign io_control_reset = reset;
  assign io_control_io_icache_read_req_valid = core_io_icache_io_read_req_valid; // @[Top.scala 19:30]
  assign io_control_io_icache_read_req_bits_addr = core_io_icache_io_read_req_bits_addr; // @[Top.scala 19:30]
  assign io_control_io_dcache_read_req_valid = core_io_dcache_io_read_req_valid; // @[Top.scala 21:30]
  assign io_control_io_dcache_read_req_bits_addr = core_io_dcache_io_read_req_bits_addr; // @[Top.scala 21:30]
  assign io_control_io_dcache_read_req_bits_rob_idx = core_io_dcache_io_read_req_bits_rob_idx; // @[Top.scala 21:30]
  assign io_control_io_dcache_write_req_valid = core_io_dcache_io_write_req_valid; // @[Top.scala 23:30]
  assign io_control_io_dcache_write_req_bits_addr = core_io_dcache_io_write_req_bits_addr; // @[Top.scala 23:30]
  assign io_control_io_dcache_write_req_bits_data = core_io_dcache_io_write_req_bits_data; // @[Top.scala 23:30]
  assign io_control_io_dcache_write_req_bits_byte_mask = core_io_dcache_io_write_req_bits_byte_mask; // @[Top.scala 23:30]
  assign io_control_io_base_ram_ctrl_data_in = io_base_ram_ctrl_data_in; // @[Top.scala 28:19]
  assign io_control_io_ext_ram_ctrl_data_in = io_ext_ram_ctrl_data_in; // @[Top.scala 27:18]
  assign io_control_io_rxd_uart_ready = io_rxd_uart_ready; // @[Top.scala 29:9]
  assign io_control_io_rxd_uart_data = io_rxd_uart_data; // @[Top.scala 29:9]
  assign io_control_io_txd_uart_busy = io_txd_uart_busy; // @[Top.scala 30:9]
  assign io_control_io_rob_commit_0_valid = core_io_rob_commit_0_valid; // @[Top.scala 25:21]
  assign io_control_io_rob_commit_0_bits_des_rob = core_io_rob_commit_0_bits_des_rob; // @[Top.scala 25:21]
  assign io_control_io_rob_commit_1_valid = core_io_rob_commit_1_valid; // @[Top.scala 25:21]
  assign io_control_io_rob_commit_1_bits_des_rob = core_io_rob_commit_1_bits_des_rob; // @[Top.scala 25:21]
  assign io_control_io_need_flush = core_io_need_flush; // @[Top.scala 24:21]
endmodule
